`timescale 1 ns/100 ps
// Version: 2022.3 2022.3.0.8


module PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM(
       W_DATA,
       R_DATA,
       W_ADDR,
       R_ADDR,
       W_EN,
       R_EN,
       CLK,
       WBYTE_EN
    );
input  [39:0] W_DATA;
output [39:0] R_DATA;
input  [15:0] W_ADDR;
input  [15:0] R_ADDR;
input  W_EN;
input  R_EN;
input  CLK;
input  [3:0] WBYTE_EN;

    wire \R_DATA_TEMPR0[0] , \R_DATA_TEMPR1[0] , \R_DATA_TEMPR2[0] , 
        \R_DATA_TEMPR3[0] , \R_DATA_TEMPR4[0] , \R_DATA_TEMPR5[0] , 
        \R_DATA_TEMPR6[0] , \R_DATA_TEMPR7[0] , \R_DATA_TEMPR8[0] , 
        \R_DATA_TEMPR9[0] , \R_DATA_TEMPR10[0] , \R_DATA_TEMPR11[0] , 
        \R_DATA_TEMPR12[0] , \R_DATA_TEMPR13[0] , \R_DATA_TEMPR14[0] , 
        \R_DATA_TEMPR15[0] , \R_DATA_TEMPR16[0] , \R_DATA_TEMPR17[0] , 
        \R_DATA_TEMPR18[0] , \R_DATA_TEMPR19[0] , \R_DATA_TEMPR20[0] , 
        \R_DATA_TEMPR21[0] , \R_DATA_TEMPR22[0] , \R_DATA_TEMPR23[0] , 
        \R_DATA_TEMPR24[0] , \R_DATA_TEMPR25[0] , \R_DATA_TEMPR26[0] , 
        \R_DATA_TEMPR27[0] , \R_DATA_TEMPR28[0] , \R_DATA_TEMPR29[0] , 
        \R_DATA_TEMPR30[0] , \R_DATA_TEMPR31[0] , \R_DATA_TEMPR32[0] , 
        \R_DATA_TEMPR33[0] , \R_DATA_TEMPR34[0] , \R_DATA_TEMPR35[0] , 
        \R_DATA_TEMPR36[0] , \R_DATA_TEMPR37[0] , \R_DATA_TEMPR38[0] , 
        \R_DATA_TEMPR39[0] , \R_DATA_TEMPR40[0] , \R_DATA_TEMPR41[0] , 
        \R_DATA_TEMPR42[0] , \R_DATA_TEMPR43[0] , \R_DATA_TEMPR44[0] , 
        \R_DATA_TEMPR45[0] , \R_DATA_TEMPR46[0] , \R_DATA_TEMPR47[0] , 
        \R_DATA_TEMPR48[0] , \R_DATA_TEMPR49[0] , \R_DATA_TEMPR50[0] , 
        \R_DATA_TEMPR51[0] , \R_DATA_TEMPR52[0] , \R_DATA_TEMPR53[0] , 
        \R_DATA_TEMPR54[0] , \R_DATA_TEMPR55[0] , \R_DATA_TEMPR56[0] , 
        \R_DATA_TEMPR57[0] , \R_DATA_TEMPR58[0] , \R_DATA_TEMPR59[0] , 
        \R_DATA_TEMPR60[0] , \R_DATA_TEMPR61[0] , \R_DATA_TEMPR62[0] , 
        \R_DATA_TEMPR63[0] , \R_DATA_TEMPR64[0] , \R_DATA_TEMPR65[0] , 
        \R_DATA_TEMPR66[0] , \R_DATA_TEMPR67[0] , \R_DATA_TEMPR68[0] , 
        \R_DATA_TEMPR69[0] , \R_DATA_TEMPR70[0] , \R_DATA_TEMPR71[0] , 
        \R_DATA_TEMPR72[0] , \R_DATA_TEMPR73[0] , \R_DATA_TEMPR74[0] , 
        \R_DATA_TEMPR75[0] , \R_DATA_TEMPR76[0] , \R_DATA_TEMPR77[0] , 
        \R_DATA_TEMPR78[0] , \R_DATA_TEMPR79[0] , \R_DATA_TEMPR80[0] , 
        \R_DATA_TEMPR81[0] , \R_DATA_TEMPR82[0] , \R_DATA_TEMPR83[0] , 
        \R_DATA_TEMPR84[0] , \R_DATA_TEMPR85[0] , \R_DATA_TEMPR86[0] , 
        \R_DATA_TEMPR87[0] , \R_DATA_TEMPR88[0] , \R_DATA_TEMPR89[0] , 
        \R_DATA_TEMPR90[0] , \R_DATA_TEMPR91[0] , \R_DATA_TEMPR92[0] , 
        \R_DATA_TEMPR93[0] , \R_DATA_TEMPR94[0] , \R_DATA_TEMPR95[0] , 
        \R_DATA_TEMPR96[0] , \R_DATA_TEMPR97[0] , \R_DATA_TEMPR98[0] , 
        \R_DATA_TEMPR99[0] , \R_DATA_TEMPR100[0] , 
        \R_DATA_TEMPR101[0] , \R_DATA_TEMPR102[0] , 
        \R_DATA_TEMPR103[0] , \R_DATA_TEMPR104[0] , 
        \R_DATA_TEMPR105[0] , \R_DATA_TEMPR106[0] , 
        \R_DATA_TEMPR107[0] , \R_DATA_TEMPR108[0] , 
        \R_DATA_TEMPR109[0] , \R_DATA_TEMPR110[0] , 
        \R_DATA_TEMPR111[0] , \R_DATA_TEMPR112[0] , 
        \R_DATA_TEMPR113[0] , \R_DATA_TEMPR114[0] , 
        \R_DATA_TEMPR115[0] , \R_DATA_TEMPR116[0] , 
        \R_DATA_TEMPR117[0] , \R_DATA_TEMPR118[0] , 
        \R_DATA_TEMPR119[0] , \R_DATA_TEMPR120[0] , 
        \R_DATA_TEMPR121[0] , \R_DATA_TEMPR122[0] , 
        \R_DATA_TEMPR123[0] , \R_DATA_TEMPR124[0] , 
        \R_DATA_TEMPR125[0] , \R_DATA_TEMPR126[0] , 
        \R_DATA_TEMPR127[0] , \R_DATA_TEMPR0[1] , \R_DATA_TEMPR1[1] , 
        \R_DATA_TEMPR2[1] , \R_DATA_TEMPR3[1] , \R_DATA_TEMPR4[1] , 
        \R_DATA_TEMPR5[1] , \R_DATA_TEMPR6[1] , \R_DATA_TEMPR7[1] , 
        \R_DATA_TEMPR8[1] , \R_DATA_TEMPR9[1] , \R_DATA_TEMPR10[1] , 
        \R_DATA_TEMPR11[1] , \R_DATA_TEMPR12[1] , \R_DATA_TEMPR13[1] , 
        \R_DATA_TEMPR14[1] , \R_DATA_TEMPR15[1] , \R_DATA_TEMPR16[1] , 
        \R_DATA_TEMPR17[1] , \R_DATA_TEMPR18[1] , \R_DATA_TEMPR19[1] , 
        \R_DATA_TEMPR20[1] , \R_DATA_TEMPR21[1] , \R_DATA_TEMPR22[1] , 
        \R_DATA_TEMPR23[1] , \R_DATA_TEMPR24[1] , \R_DATA_TEMPR25[1] , 
        \R_DATA_TEMPR26[1] , \R_DATA_TEMPR27[1] , \R_DATA_TEMPR28[1] , 
        \R_DATA_TEMPR29[1] , \R_DATA_TEMPR30[1] , \R_DATA_TEMPR31[1] , 
        \R_DATA_TEMPR32[1] , \R_DATA_TEMPR33[1] , \R_DATA_TEMPR34[1] , 
        \R_DATA_TEMPR35[1] , \R_DATA_TEMPR36[1] , \R_DATA_TEMPR37[1] , 
        \R_DATA_TEMPR38[1] , \R_DATA_TEMPR39[1] , \R_DATA_TEMPR40[1] , 
        \R_DATA_TEMPR41[1] , \R_DATA_TEMPR42[1] , \R_DATA_TEMPR43[1] , 
        \R_DATA_TEMPR44[1] , \R_DATA_TEMPR45[1] , \R_DATA_TEMPR46[1] , 
        \R_DATA_TEMPR47[1] , \R_DATA_TEMPR48[1] , \R_DATA_TEMPR49[1] , 
        \R_DATA_TEMPR50[1] , \R_DATA_TEMPR51[1] , \R_DATA_TEMPR52[1] , 
        \R_DATA_TEMPR53[1] , \R_DATA_TEMPR54[1] , \R_DATA_TEMPR55[1] , 
        \R_DATA_TEMPR56[1] , \R_DATA_TEMPR57[1] , \R_DATA_TEMPR58[1] , 
        \R_DATA_TEMPR59[1] , \R_DATA_TEMPR60[1] , \R_DATA_TEMPR61[1] , 
        \R_DATA_TEMPR62[1] , \R_DATA_TEMPR63[1] , \R_DATA_TEMPR64[1] , 
        \R_DATA_TEMPR65[1] , \R_DATA_TEMPR66[1] , \R_DATA_TEMPR67[1] , 
        \R_DATA_TEMPR68[1] , \R_DATA_TEMPR69[1] , \R_DATA_TEMPR70[1] , 
        \R_DATA_TEMPR71[1] , \R_DATA_TEMPR72[1] , \R_DATA_TEMPR73[1] , 
        \R_DATA_TEMPR74[1] , \R_DATA_TEMPR75[1] , \R_DATA_TEMPR76[1] , 
        \R_DATA_TEMPR77[1] , \R_DATA_TEMPR78[1] , \R_DATA_TEMPR79[1] , 
        \R_DATA_TEMPR80[1] , \R_DATA_TEMPR81[1] , \R_DATA_TEMPR82[1] , 
        \R_DATA_TEMPR83[1] , \R_DATA_TEMPR84[1] , \R_DATA_TEMPR85[1] , 
        \R_DATA_TEMPR86[1] , \R_DATA_TEMPR87[1] , \R_DATA_TEMPR88[1] , 
        \R_DATA_TEMPR89[1] , \R_DATA_TEMPR90[1] , \R_DATA_TEMPR91[1] , 
        \R_DATA_TEMPR92[1] , \R_DATA_TEMPR93[1] , \R_DATA_TEMPR94[1] , 
        \R_DATA_TEMPR95[1] , \R_DATA_TEMPR96[1] , \R_DATA_TEMPR97[1] , 
        \R_DATA_TEMPR98[1] , \R_DATA_TEMPR99[1] , \R_DATA_TEMPR100[1] , 
        \R_DATA_TEMPR101[1] , \R_DATA_TEMPR102[1] , 
        \R_DATA_TEMPR103[1] , \R_DATA_TEMPR104[1] , 
        \R_DATA_TEMPR105[1] , \R_DATA_TEMPR106[1] , 
        \R_DATA_TEMPR107[1] , \R_DATA_TEMPR108[1] , 
        \R_DATA_TEMPR109[1] , \R_DATA_TEMPR110[1] , 
        \R_DATA_TEMPR111[1] , \R_DATA_TEMPR112[1] , 
        \R_DATA_TEMPR113[1] , \R_DATA_TEMPR114[1] , 
        \R_DATA_TEMPR115[1] , \R_DATA_TEMPR116[1] , 
        \R_DATA_TEMPR117[1] , \R_DATA_TEMPR118[1] , 
        \R_DATA_TEMPR119[1] , \R_DATA_TEMPR120[1] , 
        \R_DATA_TEMPR121[1] , \R_DATA_TEMPR122[1] , 
        \R_DATA_TEMPR123[1] , \R_DATA_TEMPR124[1] , 
        \R_DATA_TEMPR125[1] , \R_DATA_TEMPR126[1] , 
        \R_DATA_TEMPR127[1] , \R_DATA_TEMPR0[2] , \R_DATA_TEMPR1[2] , 
        \R_DATA_TEMPR2[2] , \R_DATA_TEMPR3[2] , \R_DATA_TEMPR4[2] , 
        \R_DATA_TEMPR5[2] , \R_DATA_TEMPR6[2] , \R_DATA_TEMPR7[2] , 
        \R_DATA_TEMPR8[2] , \R_DATA_TEMPR9[2] , \R_DATA_TEMPR10[2] , 
        \R_DATA_TEMPR11[2] , \R_DATA_TEMPR12[2] , \R_DATA_TEMPR13[2] , 
        \R_DATA_TEMPR14[2] , \R_DATA_TEMPR15[2] , \R_DATA_TEMPR16[2] , 
        \R_DATA_TEMPR17[2] , \R_DATA_TEMPR18[2] , \R_DATA_TEMPR19[2] , 
        \R_DATA_TEMPR20[2] , \R_DATA_TEMPR21[2] , \R_DATA_TEMPR22[2] , 
        \R_DATA_TEMPR23[2] , \R_DATA_TEMPR24[2] , \R_DATA_TEMPR25[2] , 
        \R_DATA_TEMPR26[2] , \R_DATA_TEMPR27[2] , \R_DATA_TEMPR28[2] , 
        \R_DATA_TEMPR29[2] , \R_DATA_TEMPR30[2] , \R_DATA_TEMPR31[2] , 
        \R_DATA_TEMPR32[2] , \R_DATA_TEMPR33[2] , \R_DATA_TEMPR34[2] , 
        \R_DATA_TEMPR35[2] , \R_DATA_TEMPR36[2] , \R_DATA_TEMPR37[2] , 
        \R_DATA_TEMPR38[2] , \R_DATA_TEMPR39[2] , \R_DATA_TEMPR40[2] , 
        \R_DATA_TEMPR41[2] , \R_DATA_TEMPR42[2] , \R_DATA_TEMPR43[2] , 
        \R_DATA_TEMPR44[2] , \R_DATA_TEMPR45[2] , \R_DATA_TEMPR46[2] , 
        \R_DATA_TEMPR47[2] , \R_DATA_TEMPR48[2] , \R_DATA_TEMPR49[2] , 
        \R_DATA_TEMPR50[2] , \R_DATA_TEMPR51[2] , \R_DATA_TEMPR52[2] , 
        \R_DATA_TEMPR53[2] , \R_DATA_TEMPR54[2] , \R_DATA_TEMPR55[2] , 
        \R_DATA_TEMPR56[2] , \R_DATA_TEMPR57[2] , \R_DATA_TEMPR58[2] , 
        \R_DATA_TEMPR59[2] , \R_DATA_TEMPR60[2] , \R_DATA_TEMPR61[2] , 
        \R_DATA_TEMPR62[2] , \R_DATA_TEMPR63[2] , \R_DATA_TEMPR64[2] , 
        \R_DATA_TEMPR65[2] , \R_DATA_TEMPR66[2] , \R_DATA_TEMPR67[2] , 
        \R_DATA_TEMPR68[2] , \R_DATA_TEMPR69[2] , \R_DATA_TEMPR70[2] , 
        \R_DATA_TEMPR71[2] , \R_DATA_TEMPR72[2] , \R_DATA_TEMPR73[2] , 
        \R_DATA_TEMPR74[2] , \R_DATA_TEMPR75[2] , \R_DATA_TEMPR76[2] , 
        \R_DATA_TEMPR77[2] , \R_DATA_TEMPR78[2] , \R_DATA_TEMPR79[2] , 
        \R_DATA_TEMPR80[2] , \R_DATA_TEMPR81[2] , \R_DATA_TEMPR82[2] , 
        \R_DATA_TEMPR83[2] , \R_DATA_TEMPR84[2] , \R_DATA_TEMPR85[2] , 
        \R_DATA_TEMPR86[2] , \R_DATA_TEMPR87[2] , \R_DATA_TEMPR88[2] , 
        \R_DATA_TEMPR89[2] , \R_DATA_TEMPR90[2] , \R_DATA_TEMPR91[2] , 
        \R_DATA_TEMPR92[2] , \R_DATA_TEMPR93[2] , \R_DATA_TEMPR94[2] , 
        \R_DATA_TEMPR95[2] , \R_DATA_TEMPR96[2] , \R_DATA_TEMPR97[2] , 
        \R_DATA_TEMPR98[2] , \R_DATA_TEMPR99[2] , \R_DATA_TEMPR100[2] , 
        \R_DATA_TEMPR101[2] , \R_DATA_TEMPR102[2] , 
        \R_DATA_TEMPR103[2] , \R_DATA_TEMPR104[2] , 
        \R_DATA_TEMPR105[2] , \R_DATA_TEMPR106[2] , 
        \R_DATA_TEMPR107[2] , \R_DATA_TEMPR108[2] , 
        \R_DATA_TEMPR109[2] , \R_DATA_TEMPR110[2] , 
        \R_DATA_TEMPR111[2] , \R_DATA_TEMPR112[2] , 
        \R_DATA_TEMPR113[2] , \R_DATA_TEMPR114[2] , 
        \R_DATA_TEMPR115[2] , \R_DATA_TEMPR116[2] , 
        \R_DATA_TEMPR117[2] , \R_DATA_TEMPR118[2] , 
        \R_DATA_TEMPR119[2] , \R_DATA_TEMPR120[2] , 
        \R_DATA_TEMPR121[2] , \R_DATA_TEMPR122[2] , 
        \R_DATA_TEMPR123[2] , \R_DATA_TEMPR124[2] , 
        \R_DATA_TEMPR125[2] , \R_DATA_TEMPR126[2] , 
        \R_DATA_TEMPR127[2] , \R_DATA_TEMPR0[3] , \R_DATA_TEMPR1[3] , 
        \R_DATA_TEMPR2[3] , \R_DATA_TEMPR3[3] , \R_DATA_TEMPR4[3] , 
        \R_DATA_TEMPR5[3] , \R_DATA_TEMPR6[3] , \R_DATA_TEMPR7[3] , 
        \R_DATA_TEMPR8[3] , \R_DATA_TEMPR9[3] , \R_DATA_TEMPR10[3] , 
        \R_DATA_TEMPR11[3] , \R_DATA_TEMPR12[3] , \R_DATA_TEMPR13[3] , 
        \R_DATA_TEMPR14[3] , \R_DATA_TEMPR15[3] , \R_DATA_TEMPR16[3] , 
        \R_DATA_TEMPR17[3] , \R_DATA_TEMPR18[3] , \R_DATA_TEMPR19[3] , 
        \R_DATA_TEMPR20[3] , \R_DATA_TEMPR21[3] , \R_DATA_TEMPR22[3] , 
        \R_DATA_TEMPR23[3] , \R_DATA_TEMPR24[3] , \R_DATA_TEMPR25[3] , 
        \R_DATA_TEMPR26[3] , \R_DATA_TEMPR27[3] , \R_DATA_TEMPR28[3] , 
        \R_DATA_TEMPR29[3] , \R_DATA_TEMPR30[3] , \R_DATA_TEMPR31[3] , 
        \R_DATA_TEMPR32[3] , \R_DATA_TEMPR33[3] , \R_DATA_TEMPR34[3] , 
        \R_DATA_TEMPR35[3] , \R_DATA_TEMPR36[3] , \R_DATA_TEMPR37[3] , 
        \R_DATA_TEMPR38[3] , \R_DATA_TEMPR39[3] , \R_DATA_TEMPR40[3] , 
        \R_DATA_TEMPR41[3] , \R_DATA_TEMPR42[3] , \R_DATA_TEMPR43[3] , 
        \R_DATA_TEMPR44[3] , \R_DATA_TEMPR45[3] , \R_DATA_TEMPR46[3] , 
        \R_DATA_TEMPR47[3] , \R_DATA_TEMPR48[3] , \R_DATA_TEMPR49[3] , 
        \R_DATA_TEMPR50[3] , \R_DATA_TEMPR51[3] , \R_DATA_TEMPR52[3] , 
        \R_DATA_TEMPR53[3] , \R_DATA_TEMPR54[3] , \R_DATA_TEMPR55[3] , 
        \R_DATA_TEMPR56[3] , \R_DATA_TEMPR57[3] , \R_DATA_TEMPR58[3] , 
        \R_DATA_TEMPR59[3] , \R_DATA_TEMPR60[3] , \R_DATA_TEMPR61[3] , 
        \R_DATA_TEMPR62[3] , \R_DATA_TEMPR63[3] , \R_DATA_TEMPR64[3] , 
        \R_DATA_TEMPR65[3] , \R_DATA_TEMPR66[3] , \R_DATA_TEMPR67[3] , 
        \R_DATA_TEMPR68[3] , \R_DATA_TEMPR69[3] , \R_DATA_TEMPR70[3] , 
        \R_DATA_TEMPR71[3] , \R_DATA_TEMPR72[3] , \R_DATA_TEMPR73[3] , 
        \R_DATA_TEMPR74[3] , \R_DATA_TEMPR75[3] , \R_DATA_TEMPR76[3] , 
        \R_DATA_TEMPR77[3] , \R_DATA_TEMPR78[3] , \R_DATA_TEMPR79[3] , 
        \R_DATA_TEMPR80[3] , \R_DATA_TEMPR81[3] , \R_DATA_TEMPR82[3] , 
        \R_DATA_TEMPR83[3] , \R_DATA_TEMPR84[3] , \R_DATA_TEMPR85[3] , 
        \R_DATA_TEMPR86[3] , \R_DATA_TEMPR87[3] , \R_DATA_TEMPR88[3] , 
        \R_DATA_TEMPR89[3] , \R_DATA_TEMPR90[3] , \R_DATA_TEMPR91[3] , 
        \R_DATA_TEMPR92[3] , \R_DATA_TEMPR93[3] , \R_DATA_TEMPR94[3] , 
        \R_DATA_TEMPR95[3] , \R_DATA_TEMPR96[3] , \R_DATA_TEMPR97[3] , 
        \R_DATA_TEMPR98[3] , \R_DATA_TEMPR99[3] , \R_DATA_TEMPR100[3] , 
        \R_DATA_TEMPR101[3] , \R_DATA_TEMPR102[3] , 
        \R_DATA_TEMPR103[3] , \R_DATA_TEMPR104[3] , 
        \R_DATA_TEMPR105[3] , \R_DATA_TEMPR106[3] , 
        \R_DATA_TEMPR107[3] , \R_DATA_TEMPR108[3] , 
        \R_DATA_TEMPR109[3] , \R_DATA_TEMPR110[3] , 
        \R_DATA_TEMPR111[3] , \R_DATA_TEMPR112[3] , 
        \R_DATA_TEMPR113[3] , \R_DATA_TEMPR114[3] , 
        \R_DATA_TEMPR115[3] , \R_DATA_TEMPR116[3] , 
        \R_DATA_TEMPR117[3] , \R_DATA_TEMPR118[3] , 
        \R_DATA_TEMPR119[3] , \R_DATA_TEMPR120[3] , 
        \R_DATA_TEMPR121[3] , \R_DATA_TEMPR122[3] , 
        \R_DATA_TEMPR123[3] , \R_DATA_TEMPR124[3] , 
        \R_DATA_TEMPR125[3] , \R_DATA_TEMPR126[3] , 
        \R_DATA_TEMPR127[3] , \R_DATA_TEMPR0[4] , \R_DATA_TEMPR1[4] , 
        \R_DATA_TEMPR2[4] , \R_DATA_TEMPR3[4] , \R_DATA_TEMPR4[4] , 
        \R_DATA_TEMPR5[4] , \R_DATA_TEMPR6[4] , \R_DATA_TEMPR7[4] , 
        \R_DATA_TEMPR8[4] , \R_DATA_TEMPR9[4] , \R_DATA_TEMPR10[4] , 
        \R_DATA_TEMPR11[4] , \R_DATA_TEMPR12[4] , \R_DATA_TEMPR13[4] , 
        \R_DATA_TEMPR14[4] , \R_DATA_TEMPR15[4] , \R_DATA_TEMPR16[4] , 
        \R_DATA_TEMPR17[4] , \R_DATA_TEMPR18[4] , \R_DATA_TEMPR19[4] , 
        \R_DATA_TEMPR20[4] , \R_DATA_TEMPR21[4] , \R_DATA_TEMPR22[4] , 
        \R_DATA_TEMPR23[4] , \R_DATA_TEMPR24[4] , \R_DATA_TEMPR25[4] , 
        \R_DATA_TEMPR26[4] , \R_DATA_TEMPR27[4] , \R_DATA_TEMPR28[4] , 
        \R_DATA_TEMPR29[4] , \R_DATA_TEMPR30[4] , \R_DATA_TEMPR31[4] , 
        \R_DATA_TEMPR32[4] , \R_DATA_TEMPR33[4] , \R_DATA_TEMPR34[4] , 
        \R_DATA_TEMPR35[4] , \R_DATA_TEMPR36[4] , \R_DATA_TEMPR37[4] , 
        \R_DATA_TEMPR38[4] , \R_DATA_TEMPR39[4] , \R_DATA_TEMPR40[4] , 
        \R_DATA_TEMPR41[4] , \R_DATA_TEMPR42[4] , \R_DATA_TEMPR43[4] , 
        \R_DATA_TEMPR44[4] , \R_DATA_TEMPR45[4] , \R_DATA_TEMPR46[4] , 
        \R_DATA_TEMPR47[4] , \R_DATA_TEMPR48[4] , \R_DATA_TEMPR49[4] , 
        \R_DATA_TEMPR50[4] , \R_DATA_TEMPR51[4] , \R_DATA_TEMPR52[4] , 
        \R_DATA_TEMPR53[4] , \R_DATA_TEMPR54[4] , \R_DATA_TEMPR55[4] , 
        \R_DATA_TEMPR56[4] , \R_DATA_TEMPR57[4] , \R_DATA_TEMPR58[4] , 
        \R_DATA_TEMPR59[4] , \R_DATA_TEMPR60[4] , \R_DATA_TEMPR61[4] , 
        \R_DATA_TEMPR62[4] , \R_DATA_TEMPR63[4] , \R_DATA_TEMPR64[4] , 
        \R_DATA_TEMPR65[4] , \R_DATA_TEMPR66[4] , \R_DATA_TEMPR67[4] , 
        \R_DATA_TEMPR68[4] , \R_DATA_TEMPR69[4] , \R_DATA_TEMPR70[4] , 
        \R_DATA_TEMPR71[4] , \R_DATA_TEMPR72[4] , \R_DATA_TEMPR73[4] , 
        \R_DATA_TEMPR74[4] , \R_DATA_TEMPR75[4] , \R_DATA_TEMPR76[4] , 
        \R_DATA_TEMPR77[4] , \R_DATA_TEMPR78[4] , \R_DATA_TEMPR79[4] , 
        \R_DATA_TEMPR80[4] , \R_DATA_TEMPR81[4] , \R_DATA_TEMPR82[4] , 
        \R_DATA_TEMPR83[4] , \R_DATA_TEMPR84[4] , \R_DATA_TEMPR85[4] , 
        \R_DATA_TEMPR86[4] , \R_DATA_TEMPR87[4] , \R_DATA_TEMPR88[4] , 
        \R_DATA_TEMPR89[4] , \R_DATA_TEMPR90[4] , \R_DATA_TEMPR91[4] , 
        \R_DATA_TEMPR92[4] , \R_DATA_TEMPR93[4] , \R_DATA_TEMPR94[4] , 
        \R_DATA_TEMPR95[4] , \R_DATA_TEMPR96[4] , \R_DATA_TEMPR97[4] , 
        \R_DATA_TEMPR98[4] , \R_DATA_TEMPR99[4] , \R_DATA_TEMPR100[4] , 
        \R_DATA_TEMPR101[4] , \R_DATA_TEMPR102[4] , 
        \R_DATA_TEMPR103[4] , \R_DATA_TEMPR104[4] , 
        \R_DATA_TEMPR105[4] , \R_DATA_TEMPR106[4] , 
        \R_DATA_TEMPR107[4] , \R_DATA_TEMPR108[4] , 
        \R_DATA_TEMPR109[4] , \R_DATA_TEMPR110[4] , 
        \R_DATA_TEMPR111[4] , \R_DATA_TEMPR112[4] , 
        \R_DATA_TEMPR113[4] , \R_DATA_TEMPR114[4] , 
        \R_DATA_TEMPR115[4] , \R_DATA_TEMPR116[4] , 
        \R_DATA_TEMPR117[4] , \R_DATA_TEMPR118[4] , 
        \R_DATA_TEMPR119[4] , \R_DATA_TEMPR120[4] , 
        \R_DATA_TEMPR121[4] , \R_DATA_TEMPR122[4] , 
        \R_DATA_TEMPR123[4] , \R_DATA_TEMPR124[4] , 
        \R_DATA_TEMPR125[4] , \R_DATA_TEMPR126[4] , 
        \R_DATA_TEMPR127[4] , \R_DATA_TEMPR0[5] , \R_DATA_TEMPR1[5] , 
        \R_DATA_TEMPR2[5] , \R_DATA_TEMPR3[5] , \R_DATA_TEMPR4[5] , 
        \R_DATA_TEMPR5[5] , \R_DATA_TEMPR6[5] , \R_DATA_TEMPR7[5] , 
        \R_DATA_TEMPR8[5] , \R_DATA_TEMPR9[5] , \R_DATA_TEMPR10[5] , 
        \R_DATA_TEMPR11[5] , \R_DATA_TEMPR12[5] , \R_DATA_TEMPR13[5] , 
        \R_DATA_TEMPR14[5] , \R_DATA_TEMPR15[5] , \R_DATA_TEMPR16[5] , 
        \R_DATA_TEMPR17[5] , \R_DATA_TEMPR18[5] , \R_DATA_TEMPR19[5] , 
        \R_DATA_TEMPR20[5] , \R_DATA_TEMPR21[5] , \R_DATA_TEMPR22[5] , 
        \R_DATA_TEMPR23[5] , \R_DATA_TEMPR24[5] , \R_DATA_TEMPR25[5] , 
        \R_DATA_TEMPR26[5] , \R_DATA_TEMPR27[5] , \R_DATA_TEMPR28[5] , 
        \R_DATA_TEMPR29[5] , \R_DATA_TEMPR30[5] , \R_DATA_TEMPR31[5] , 
        \R_DATA_TEMPR32[5] , \R_DATA_TEMPR33[5] , \R_DATA_TEMPR34[5] , 
        \R_DATA_TEMPR35[5] , \R_DATA_TEMPR36[5] , \R_DATA_TEMPR37[5] , 
        \R_DATA_TEMPR38[5] , \R_DATA_TEMPR39[5] , \R_DATA_TEMPR40[5] , 
        \R_DATA_TEMPR41[5] , \R_DATA_TEMPR42[5] , \R_DATA_TEMPR43[5] , 
        \R_DATA_TEMPR44[5] , \R_DATA_TEMPR45[5] , \R_DATA_TEMPR46[5] , 
        \R_DATA_TEMPR47[5] , \R_DATA_TEMPR48[5] , \R_DATA_TEMPR49[5] , 
        \R_DATA_TEMPR50[5] , \R_DATA_TEMPR51[5] , \R_DATA_TEMPR52[5] , 
        \R_DATA_TEMPR53[5] , \R_DATA_TEMPR54[5] , \R_DATA_TEMPR55[5] , 
        \R_DATA_TEMPR56[5] , \R_DATA_TEMPR57[5] , \R_DATA_TEMPR58[5] , 
        \R_DATA_TEMPR59[5] , \R_DATA_TEMPR60[5] , \R_DATA_TEMPR61[5] , 
        \R_DATA_TEMPR62[5] , \R_DATA_TEMPR63[5] , \R_DATA_TEMPR64[5] , 
        \R_DATA_TEMPR65[5] , \R_DATA_TEMPR66[5] , \R_DATA_TEMPR67[5] , 
        \R_DATA_TEMPR68[5] , \R_DATA_TEMPR69[5] , \R_DATA_TEMPR70[5] , 
        \R_DATA_TEMPR71[5] , \R_DATA_TEMPR72[5] , \R_DATA_TEMPR73[5] , 
        \R_DATA_TEMPR74[5] , \R_DATA_TEMPR75[5] , \R_DATA_TEMPR76[5] , 
        \R_DATA_TEMPR77[5] , \R_DATA_TEMPR78[5] , \R_DATA_TEMPR79[5] , 
        \R_DATA_TEMPR80[5] , \R_DATA_TEMPR81[5] , \R_DATA_TEMPR82[5] , 
        \R_DATA_TEMPR83[5] , \R_DATA_TEMPR84[5] , \R_DATA_TEMPR85[5] , 
        \R_DATA_TEMPR86[5] , \R_DATA_TEMPR87[5] , \R_DATA_TEMPR88[5] , 
        \R_DATA_TEMPR89[5] , \R_DATA_TEMPR90[5] , \R_DATA_TEMPR91[5] , 
        \R_DATA_TEMPR92[5] , \R_DATA_TEMPR93[5] , \R_DATA_TEMPR94[5] , 
        \R_DATA_TEMPR95[5] , \R_DATA_TEMPR96[5] , \R_DATA_TEMPR97[5] , 
        \R_DATA_TEMPR98[5] , \R_DATA_TEMPR99[5] , \R_DATA_TEMPR100[5] , 
        \R_DATA_TEMPR101[5] , \R_DATA_TEMPR102[5] , 
        \R_DATA_TEMPR103[5] , \R_DATA_TEMPR104[5] , 
        \R_DATA_TEMPR105[5] , \R_DATA_TEMPR106[5] , 
        \R_DATA_TEMPR107[5] , \R_DATA_TEMPR108[5] , 
        \R_DATA_TEMPR109[5] , \R_DATA_TEMPR110[5] , 
        \R_DATA_TEMPR111[5] , \R_DATA_TEMPR112[5] , 
        \R_DATA_TEMPR113[5] , \R_DATA_TEMPR114[5] , 
        \R_DATA_TEMPR115[5] , \R_DATA_TEMPR116[5] , 
        \R_DATA_TEMPR117[5] , \R_DATA_TEMPR118[5] , 
        \R_DATA_TEMPR119[5] , \R_DATA_TEMPR120[5] , 
        \R_DATA_TEMPR121[5] , \R_DATA_TEMPR122[5] , 
        \R_DATA_TEMPR123[5] , \R_DATA_TEMPR124[5] , 
        \R_DATA_TEMPR125[5] , \R_DATA_TEMPR126[5] , 
        \R_DATA_TEMPR127[5] , \R_DATA_TEMPR0[6] , \R_DATA_TEMPR1[6] , 
        \R_DATA_TEMPR2[6] , \R_DATA_TEMPR3[6] , \R_DATA_TEMPR4[6] , 
        \R_DATA_TEMPR5[6] , \R_DATA_TEMPR6[6] , \R_DATA_TEMPR7[6] , 
        \R_DATA_TEMPR8[6] , \R_DATA_TEMPR9[6] , \R_DATA_TEMPR10[6] , 
        \R_DATA_TEMPR11[6] , \R_DATA_TEMPR12[6] , \R_DATA_TEMPR13[6] , 
        \R_DATA_TEMPR14[6] , \R_DATA_TEMPR15[6] , \R_DATA_TEMPR16[6] , 
        \R_DATA_TEMPR17[6] , \R_DATA_TEMPR18[6] , \R_DATA_TEMPR19[6] , 
        \R_DATA_TEMPR20[6] , \R_DATA_TEMPR21[6] , \R_DATA_TEMPR22[6] , 
        \R_DATA_TEMPR23[6] , \R_DATA_TEMPR24[6] , \R_DATA_TEMPR25[6] , 
        \R_DATA_TEMPR26[6] , \R_DATA_TEMPR27[6] , \R_DATA_TEMPR28[6] , 
        \R_DATA_TEMPR29[6] , \R_DATA_TEMPR30[6] , \R_DATA_TEMPR31[6] , 
        \R_DATA_TEMPR32[6] , \R_DATA_TEMPR33[6] , \R_DATA_TEMPR34[6] , 
        \R_DATA_TEMPR35[6] , \R_DATA_TEMPR36[6] , \R_DATA_TEMPR37[6] , 
        \R_DATA_TEMPR38[6] , \R_DATA_TEMPR39[6] , \R_DATA_TEMPR40[6] , 
        \R_DATA_TEMPR41[6] , \R_DATA_TEMPR42[6] , \R_DATA_TEMPR43[6] , 
        \R_DATA_TEMPR44[6] , \R_DATA_TEMPR45[6] , \R_DATA_TEMPR46[6] , 
        \R_DATA_TEMPR47[6] , \R_DATA_TEMPR48[6] , \R_DATA_TEMPR49[6] , 
        \R_DATA_TEMPR50[6] , \R_DATA_TEMPR51[6] , \R_DATA_TEMPR52[6] , 
        \R_DATA_TEMPR53[6] , \R_DATA_TEMPR54[6] , \R_DATA_TEMPR55[6] , 
        \R_DATA_TEMPR56[6] , \R_DATA_TEMPR57[6] , \R_DATA_TEMPR58[6] , 
        \R_DATA_TEMPR59[6] , \R_DATA_TEMPR60[6] , \R_DATA_TEMPR61[6] , 
        \R_DATA_TEMPR62[6] , \R_DATA_TEMPR63[6] , \R_DATA_TEMPR64[6] , 
        \R_DATA_TEMPR65[6] , \R_DATA_TEMPR66[6] , \R_DATA_TEMPR67[6] , 
        \R_DATA_TEMPR68[6] , \R_DATA_TEMPR69[6] , \R_DATA_TEMPR70[6] , 
        \R_DATA_TEMPR71[6] , \R_DATA_TEMPR72[6] , \R_DATA_TEMPR73[6] , 
        \R_DATA_TEMPR74[6] , \R_DATA_TEMPR75[6] , \R_DATA_TEMPR76[6] , 
        \R_DATA_TEMPR77[6] , \R_DATA_TEMPR78[6] , \R_DATA_TEMPR79[6] , 
        \R_DATA_TEMPR80[6] , \R_DATA_TEMPR81[6] , \R_DATA_TEMPR82[6] , 
        \R_DATA_TEMPR83[6] , \R_DATA_TEMPR84[6] , \R_DATA_TEMPR85[6] , 
        \R_DATA_TEMPR86[6] , \R_DATA_TEMPR87[6] , \R_DATA_TEMPR88[6] , 
        \R_DATA_TEMPR89[6] , \R_DATA_TEMPR90[6] , \R_DATA_TEMPR91[6] , 
        \R_DATA_TEMPR92[6] , \R_DATA_TEMPR93[6] , \R_DATA_TEMPR94[6] , 
        \R_DATA_TEMPR95[6] , \R_DATA_TEMPR96[6] , \R_DATA_TEMPR97[6] , 
        \R_DATA_TEMPR98[6] , \R_DATA_TEMPR99[6] , \R_DATA_TEMPR100[6] , 
        \R_DATA_TEMPR101[6] , \R_DATA_TEMPR102[6] , 
        \R_DATA_TEMPR103[6] , \R_DATA_TEMPR104[6] , 
        \R_DATA_TEMPR105[6] , \R_DATA_TEMPR106[6] , 
        \R_DATA_TEMPR107[6] , \R_DATA_TEMPR108[6] , 
        \R_DATA_TEMPR109[6] , \R_DATA_TEMPR110[6] , 
        \R_DATA_TEMPR111[6] , \R_DATA_TEMPR112[6] , 
        \R_DATA_TEMPR113[6] , \R_DATA_TEMPR114[6] , 
        \R_DATA_TEMPR115[6] , \R_DATA_TEMPR116[6] , 
        \R_DATA_TEMPR117[6] , \R_DATA_TEMPR118[6] , 
        \R_DATA_TEMPR119[6] , \R_DATA_TEMPR120[6] , 
        \R_DATA_TEMPR121[6] , \R_DATA_TEMPR122[6] , 
        \R_DATA_TEMPR123[6] , \R_DATA_TEMPR124[6] , 
        \R_DATA_TEMPR125[6] , \R_DATA_TEMPR126[6] , 
        \R_DATA_TEMPR127[6] , \R_DATA_TEMPR0[7] , \R_DATA_TEMPR1[7] , 
        \R_DATA_TEMPR2[7] , \R_DATA_TEMPR3[7] , \R_DATA_TEMPR4[7] , 
        \R_DATA_TEMPR5[7] , \R_DATA_TEMPR6[7] , \R_DATA_TEMPR7[7] , 
        \R_DATA_TEMPR8[7] , \R_DATA_TEMPR9[7] , \R_DATA_TEMPR10[7] , 
        \R_DATA_TEMPR11[7] , \R_DATA_TEMPR12[7] , \R_DATA_TEMPR13[7] , 
        \R_DATA_TEMPR14[7] , \R_DATA_TEMPR15[7] , \R_DATA_TEMPR16[7] , 
        \R_DATA_TEMPR17[7] , \R_DATA_TEMPR18[7] , \R_DATA_TEMPR19[7] , 
        \R_DATA_TEMPR20[7] , \R_DATA_TEMPR21[7] , \R_DATA_TEMPR22[7] , 
        \R_DATA_TEMPR23[7] , \R_DATA_TEMPR24[7] , \R_DATA_TEMPR25[7] , 
        \R_DATA_TEMPR26[7] , \R_DATA_TEMPR27[7] , \R_DATA_TEMPR28[7] , 
        \R_DATA_TEMPR29[7] , \R_DATA_TEMPR30[7] , \R_DATA_TEMPR31[7] , 
        \R_DATA_TEMPR32[7] , \R_DATA_TEMPR33[7] , \R_DATA_TEMPR34[7] , 
        \R_DATA_TEMPR35[7] , \R_DATA_TEMPR36[7] , \R_DATA_TEMPR37[7] , 
        \R_DATA_TEMPR38[7] , \R_DATA_TEMPR39[7] , \R_DATA_TEMPR40[7] , 
        \R_DATA_TEMPR41[7] , \R_DATA_TEMPR42[7] , \R_DATA_TEMPR43[7] , 
        \R_DATA_TEMPR44[7] , \R_DATA_TEMPR45[7] , \R_DATA_TEMPR46[7] , 
        \R_DATA_TEMPR47[7] , \R_DATA_TEMPR48[7] , \R_DATA_TEMPR49[7] , 
        \R_DATA_TEMPR50[7] , \R_DATA_TEMPR51[7] , \R_DATA_TEMPR52[7] , 
        \R_DATA_TEMPR53[7] , \R_DATA_TEMPR54[7] , \R_DATA_TEMPR55[7] , 
        \R_DATA_TEMPR56[7] , \R_DATA_TEMPR57[7] , \R_DATA_TEMPR58[7] , 
        \R_DATA_TEMPR59[7] , \R_DATA_TEMPR60[7] , \R_DATA_TEMPR61[7] , 
        \R_DATA_TEMPR62[7] , \R_DATA_TEMPR63[7] , \R_DATA_TEMPR64[7] , 
        \R_DATA_TEMPR65[7] , \R_DATA_TEMPR66[7] , \R_DATA_TEMPR67[7] , 
        \R_DATA_TEMPR68[7] , \R_DATA_TEMPR69[7] , \R_DATA_TEMPR70[7] , 
        \R_DATA_TEMPR71[7] , \R_DATA_TEMPR72[7] , \R_DATA_TEMPR73[7] , 
        \R_DATA_TEMPR74[7] , \R_DATA_TEMPR75[7] , \R_DATA_TEMPR76[7] , 
        \R_DATA_TEMPR77[7] , \R_DATA_TEMPR78[7] , \R_DATA_TEMPR79[7] , 
        \R_DATA_TEMPR80[7] , \R_DATA_TEMPR81[7] , \R_DATA_TEMPR82[7] , 
        \R_DATA_TEMPR83[7] , \R_DATA_TEMPR84[7] , \R_DATA_TEMPR85[7] , 
        \R_DATA_TEMPR86[7] , \R_DATA_TEMPR87[7] , \R_DATA_TEMPR88[7] , 
        \R_DATA_TEMPR89[7] , \R_DATA_TEMPR90[7] , \R_DATA_TEMPR91[7] , 
        \R_DATA_TEMPR92[7] , \R_DATA_TEMPR93[7] , \R_DATA_TEMPR94[7] , 
        \R_DATA_TEMPR95[7] , \R_DATA_TEMPR96[7] , \R_DATA_TEMPR97[7] , 
        \R_DATA_TEMPR98[7] , \R_DATA_TEMPR99[7] , \R_DATA_TEMPR100[7] , 
        \R_DATA_TEMPR101[7] , \R_DATA_TEMPR102[7] , 
        \R_DATA_TEMPR103[7] , \R_DATA_TEMPR104[7] , 
        \R_DATA_TEMPR105[7] , \R_DATA_TEMPR106[7] , 
        \R_DATA_TEMPR107[7] , \R_DATA_TEMPR108[7] , 
        \R_DATA_TEMPR109[7] , \R_DATA_TEMPR110[7] , 
        \R_DATA_TEMPR111[7] , \R_DATA_TEMPR112[7] , 
        \R_DATA_TEMPR113[7] , \R_DATA_TEMPR114[7] , 
        \R_DATA_TEMPR115[7] , \R_DATA_TEMPR116[7] , 
        \R_DATA_TEMPR117[7] , \R_DATA_TEMPR118[7] , 
        \R_DATA_TEMPR119[7] , \R_DATA_TEMPR120[7] , 
        \R_DATA_TEMPR121[7] , \R_DATA_TEMPR122[7] , 
        \R_DATA_TEMPR123[7] , \R_DATA_TEMPR124[7] , 
        \R_DATA_TEMPR125[7] , \R_DATA_TEMPR126[7] , 
        \R_DATA_TEMPR127[7] , \R_DATA_TEMPR0[8] , \R_DATA_TEMPR1[8] , 
        \R_DATA_TEMPR2[8] , \R_DATA_TEMPR3[8] , \R_DATA_TEMPR4[8] , 
        \R_DATA_TEMPR5[8] , \R_DATA_TEMPR6[8] , \R_DATA_TEMPR7[8] , 
        \R_DATA_TEMPR8[8] , \R_DATA_TEMPR9[8] , \R_DATA_TEMPR10[8] , 
        \R_DATA_TEMPR11[8] , \R_DATA_TEMPR12[8] , \R_DATA_TEMPR13[8] , 
        \R_DATA_TEMPR14[8] , \R_DATA_TEMPR15[8] , \R_DATA_TEMPR16[8] , 
        \R_DATA_TEMPR17[8] , \R_DATA_TEMPR18[8] , \R_DATA_TEMPR19[8] , 
        \R_DATA_TEMPR20[8] , \R_DATA_TEMPR21[8] , \R_DATA_TEMPR22[8] , 
        \R_DATA_TEMPR23[8] , \R_DATA_TEMPR24[8] , \R_DATA_TEMPR25[8] , 
        \R_DATA_TEMPR26[8] , \R_DATA_TEMPR27[8] , \R_DATA_TEMPR28[8] , 
        \R_DATA_TEMPR29[8] , \R_DATA_TEMPR30[8] , \R_DATA_TEMPR31[8] , 
        \R_DATA_TEMPR32[8] , \R_DATA_TEMPR33[8] , \R_DATA_TEMPR34[8] , 
        \R_DATA_TEMPR35[8] , \R_DATA_TEMPR36[8] , \R_DATA_TEMPR37[8] , 
        \R_DATA_TEMPR38[8] , \R_DATA_TEMPR39[8] , \R_DATA_TEMPR40[8] , 
        \R_DATA_TEMPR41[8] , \R_DATA_TEMPR42[8] , \R_DATA_TEMPR43[8] , 
        \R_DATA_TEMPR44[8] , \R_DATA_TEMPR45[8] , \R_DATA_TEMPR46[8] , 
        \R_DATA_TEMPR47[8] , \R_DATA_TEMPR48[8] , \R_DATA_TEMPR49[8] , 
        \R_DATA_TEMPR50[8] , \R_DATA_TEMPR51[8] , \R_DATA_TEMPR52[8] , 
        \R_DATA_TEMPR53[8] , \R_DATA_TEMPR54[8] , \R_DATA_TEMPR55[8] , 
        \R_DATA_TEMPR56[8] , \R_DATA_TEMPR57[8] , \R_DATA_TEMPR58[8] , 
        \R_DATA_TEMPR59[8] , \R_DATA_TEMPR60[8] , \R_DATA_TEMPR61[8] , 
        \R_DATA_TEMPR62[8] , \R_DATA_TEMPR63[8] , \R_DATA_TEMPR64[8] , 
        \R_DATA_TEMPR65[8] , \R_DATA_TEMPR66[8] , \R_DATA_TEMPR67[8] , 
        \R_DATA_TEMPR68[8] , \R_DATA_TEMPR69[8] , \R_DATA_TEMPR70[8] , 
        \R_DATA_TEMPR71[8] , \R_DATA_TEMPR72[8] , \R_DATA_TEMPR73[8] , 
        \R_DATA_TEMPR74[8] , \R_DATA_TEMPR75[8] , \R_DATA_TEMPR76[8] , 
        \R_DATA_TEMPR77[8] , \R_DATA_TEMPR78[8] , \R_DATA_TEMPR79[8] , 
        \R_DATA_TEMPR80[8] , \R_DATA_TEMPR81[8] , \R_DATA_TEMPR82[8] , 
        \R_DATA_TEMPR83[8] , \R_DATA_TEMPR84[8] , \R_DATA_TEMPR85[8] , 
        \R_DATA_TEMPR86[8] , \R_DATA_TEMPR87[8] , \R_DATA_TEMPR88[8] , 
        \R_DATA_TEMPR89[8] , \R_DATA_TEMPR90[8] , \R_DATA_TEMPR91[8] , 
        \R_DATA_TEMPR92[8] , \R_DATA_TEMPR93[8] , \R_DATA_TEMPR94[8] , 
        \R_DATA_TEMPR95[8] , \R_DATA_TEMPR96[8] , \R_DATA_TEMPR97[8] , 
        \R_DATA_TEMPR98[8] , \R_DATA_TEMPR99[8] , \R_DATA_TEMPR100[8] , 
        \R_DATA_TEMPR101[8] , \R_DATA_TEMPR102[8] , 
        \R_DATA_TEMPR103[8] , \R_DATA_TEMPR104[8] , 
        \R_DATA_TEMPR105[8] , \R_DATA_TEMPR106[8] , 
        \R_DATA_TEMPR107[8] , \R_DATA_TEMPR108[8] , 
        \R_DATA_TEMPR109[8] , \R_DATA_TEMPR110[8] , 
        \R_DATA_TEMPR111[8] , \R_DATA_TEMPR112[8] , 
        \R_DATA_TEMPR113[8] , \R_DATA_TEMPR114[8] , 
        \R_DATA_TEMPR115[8] , \R_DATA_TEMPR116[8] , 
        \R_DATA_TEMPR117[8] , \R_DATA_TEMPR118[8] , 
        \R_DATA_TEMPR119[8] , \R_DATA_TEMPR120[8] , 
        \R_DATA_TEMPR121[8] , \R_DATA_TEMPR122[8] , 
        \R_DATA_TEMPR123[8] , \R_DATA_TEMPR124[8] , 
        \R_DATA_TEMPR125[8] , \R_DATA_TEMPR126[8] , 
        \R_DATA_TEMPR127[8] , \R_DATA_TEMPR0[9] , \R_DATA_TEMPR1[9] , 
        \R_DATA_TEMPR2[9] , \R_DATA_TEMPR3[9] , \R_DATA_TEMPR4[9] , 
        \R_DATA_TEMPR5[9] , \R_DATA_TEMPR6[9] , \R_DATA_TEMPR7[9] , 
        \R_DATA_TEMPR8[9] , \R_DATA_TEMPR9[9] , \R_DATA_TEMPR10[9] , 
        \R_DATA_TEMPR11[9] , \R_DATA_TEMPR12[9] , \R_DATA_TEMPR13[9] , 
        \R_DATA_TEMPR14[9] , \R_DATA_TEMPR15[9] , \R_DATA_TEMPR16[9] , 
        \R_DATA_TEMPR17[9] , \R_DATA_TEMPR18[9] , \R_DATA_TEMPR19[9] , 
        \R_DATA_TEMPR20[9] , \R_DATA_TEMPR21[9] , \R_DATA_TEMPR22[9] , 
        \R_DATA_TEMPR23[9] , \R_DATA_TEMPR24[9] , \R_DATA_TEMPR25[9] , 
        \R_DATA_TEMPR26[9] , \R_DATA_TEMPR27[9] , \R_DATA_TEMPR28[9] , 
        \R_DATA_TEMPR29[9] , \R_DATA_TEMPR30[9] , \R_DATA_TEMPR31[9] , 
        \R_DATA_TEMPR32[9] , \R_DATA_TEMPR33[9] , \R_DATA_TEMPR34[9] , 
        \R_DATA_TEMPR35[9] , \R_DATA_TEMPR36[9] , \R_DATA_TEMPR37[9] , 
        \R_DATA_TEMPR38[9] , \R_DATA_TEMPR39[9] , \R_DATA_TEMPR40[9] , 
        \R_DATA_TEMPR41[9] , \R_DATA_TEMPR42[9] , \R_DATA_TEMPR43[9] , 
        \R_DATA_TEMPR44[9] , \R_DATA_TEMPR45[9] , \R_DATA_TEMPR46[9] , 
        \R_DATA_TEMPR47[9] , \R_DATA_TEMPR48[9] , \R_DATA_TEMPR49[9] , 
        \R_DATA_TEMPR50[9] , \R_DATA_TEMPR51[9] , \R_DATA_TEMPR52[9] , 
        \R_DATA_TEMPR53[9] , \R_DATA_TEMPR54[9] , \R_DATA_TEMPR55[9] , 
        \R_DATA_TEMPR56[9] , \R_DATA_TEMPR57[9] , \R_DATA_TEMPR58[9] , 
        \R_DATA_TEMPR59[9] , \R_DATA_TEMPR60[9] , \R_DATA_TEMPR61[9] , 
        \R_DATA_TEMPR62[9] , \R_DATA_TEMPR63[9] , \R_DATA_TEMPR64[9] , 
        \R_DATA_TEMPR65[9] , \R_DATA_TEMPR66[9] , \R_DATA_TEMPR67[9] , 
        \R_DATA_TEMPR68[9] , \R_DATA_TEMPR69[9] , \R_DATA_TEMPR70[9] , 
        \R_DATA_TEMPR71[9] , \R_DATA_TEMPR72[9] , \R_DATA_TEMPR73[9] , 
        \R_DATA_TEMPR74[9] , \R_DATA_TEMPR75[9] , \R_DATA_TEMPR76[9] , 
        \R_DATA_TEMPR77[9] , \R_DATA_TEMPR78[9] , \R_DATA_TEMPR79[9] , 
        \R_DATA_TEMPR80[9] , \R_DATA_TEMPR81[9] , \R_DATA_TEMPR82[9] , 
        \R_DATA_TEMPR83[9] , \R_DATA_TEMPR84[9] , \R_DATA_TEMPR85[9] , 
        \R_DATA_TEMPR86[9] , \R_DATA_TEMPR87[9] , \R_DATA_TEMPR88[9] , 
        \R_DATA_TEMPR89[9] , \R_DATA_TEMPR90[9] , \R_DATA_TEMPR91[9] , 
        \R_DATA_TEMPR92[9] , \R_DATA_TEMPR93[9] , \R_DATA_TEMPR94[9] , 
        \R_DATA_TEMPR95[9] , \R_DATA_TEMPR96[9] , \R_DATA_TEMPR97[9] , 
        \R_DATA_TEMPR98[9] , \R_DATA_TEMPR99[9] , \R_DATA_TEMPR100[9] , 
        \R_DATA_TEMPR101[9] , \R_DATA_TEMPR102[9] , 
        \R_DATA_TEMPR103[9] , \R_DATA_TEMPR104[9] , 
        \R_DATA_TEMPR105[9] , \R_DATA_TEMPR106[9] , 
        \R_DATA_TEMPR107[9] , \R_DATA_TEMPR108[9] , 
        \R_DATA_TEMPR109[9] , \R_DATA_TEMPR110[9] , 
        \R_DATA_TEMPR111[9] , \R_DATA_TEMPR112[9] , 
        \R_DATA_TEMPR113[9] , \R_DATA_TEMPR114[9] , 
        \R_DATA_TEMPR115[9] , \R_DATA_TEMPR116[9] , 
        \R_DATA_TEMPR117[9] , \R_DATA_TEMPR118[9] , 
        \R_DATA_TEMPR119[9] , \R_DATA_TEMPR120[9] , 
        \R_DATA_TEMPR121[9] , \R_DATA_TEMPR122[9] , 
        \R_DATA_TEMPR123[9] , \R_DATA_TEMPR124[9] , 
        \R_DATA_TEMPR125[9] , \R_DATA_TEMPR126[9] , 
        \R_DATA_TEMPR127[9] , \R_DATA_TEMPR0[10] , \R_DATA_TEMPR1[10] , 
        \R_DATA_TEMPR2[10] , \R_DATA_TEMPR3[10] , \R_DATA_TEMPR4[10] , 
        \R_DATA_TEMPR5[10] , \R_DATA_TEMPR6[10] , \R_DATA_TEMPR7[10] , 
        \R_DATA_TEMPR8[10] , \R_DATA_TEMPR9[10] , \R_DATA_TEMPR10[10] , 
        \R_DATA_TEMPR11[10] , \R_DATA_TEMPR12[10] , 
        \R_DATA_TEMPR13[10] , \R_DATA_TEMPR14[10] , 
        \R_DATA_TEMPR15[10] , \R_DATA_TEMPR16[10] , 
        \R_DATA_TEMPR17[10] , \R_DATA_TEMPR18[10] , 
        \R_DATA_TEMPR19[10] , \R_DATA_TEMPR20[10] , 
        \R_DATA_TEMPR21[10] , \R_DATA_TEMPR22[10] , 
        \R_DATA_TEMPR23[10] , \R_DATA_TEMPR24[10] , 
        \R_DATA_TEMPR25[10] , \R_DATA_TEMPR26[10] , 
        \R_DATA_TEMPR27[10] , \R_DATA_TEMPR28[10] , 
        \R_DATA_TEMPR29[10] , \R_DATA_TEMPR30[10] , 
        \R_DATA_TEMPR31[10] , \R_DATA_TEMPR32[10] , 
        \R_DATA_TEMPR33[10] , \R_DATA_TEMPR34[10] , 
        \R_DATA_TEMPR35[10] , \R_DATA_TEMPR36[10] , 
        \R_DATA_TEMPR37[10] , \R_DATA_TEMPR38[10] , 
        \R_DATA_TEMPR39[10] , \R_DATA_TEMPR40[10] , 
        \R_DATA_TEMPR41[10] , \R_DATA_TEMPR42[10] , 
        \R_DATA_TEMPR43[10] , \R_DATA_TEMPR44[10] , 
        \R_DATA_TEMPR45[10] , \R_DATA_TEMPR46[10] , 
        \R_DATA_TEMPR47[10] , \R_DATA_TEMPR48[10] , 
        \R_DATA_TEMPR49[10] , \R_DATA_TEMPR50[10] , 
        \R_DATA_TEMPR51[10] , \R_DATA_TEMPR52[10] , 
        \R_DATA_TEMPR53[10] , \R_DATA_TEMPR54[10] , 
        \R_DATA_TEMPR55[10] , \R_DATA_TEMPR56[10] , 
        \R_DATA_TEMPR57[10] , \R_DATA_TEMPR58[10] , 
        \R_DATA_TEMPR59[10] , \R_DATA_TEMPR60[10] , 
        \R_DATA_TEMPR61[10] , \R_DATA_TEMPR62[10] , 
        \R_DATA_TEMPR63[10] , \R_DATA_TEMPR64[10] , 
        \R_DATA_TEMPR65[10] , \R_DATA_TEMPR66[10] , 
        \R_DATA_TEMPR67[10] , \R_DATA_TEMPR68[10] , 
        \R_DATA_TEMPR69[10] , \R_DATA_TEMPR70[10] , 
        \R_DATA_TEMPR71[10] , \R_DATA_TEMPR72[10] , 
        \R_DATA_TEMPR73[10] , \R_DATA_TEMPR74[10] , 
        \R_DATA_TEMPR75[10] , \R_DATA_TEMPR76[10] , 
        \R_DATA_TEMPR77[10] , \R_DATA_TEMPR78[10] , 
        \R_DATA_TEMPR79[10] , \R_DATA_TEMPR80[10] , 
        \R_DATA_TEMPR81[10] , \R_DATA_TEMPR82[10] , 
        \R_DATA_TEMPR83[10] , \R_DATA_TEMPR84[10] , 
        \R_DATA_TEMPR85[10] , \R_DATA_TEMPR86[10] , 
        \R_DATA_TEMPR87[10] , \R_DATA_TEMPR88[10] , 
        \R_DATA_TEMPR89[10] , \R_DATA_TEMPR90[10] , 
        \R_DATA_TEMPR91[10] , \R_DATA_TEMPR92[10] , 
        \R_DATA_TEMPR93[10] , \R_DATA_TEMPR94[10] , 
        \R_DATA_TEMPR95[10] , \R_DATA_TEMPR96[10] , 
        \R_DATA_TEMPR97[10] , \R_DATA_TEMPR98[10] , 
        \R_DATA_TEMPR99[10] , \R_DATA_TEMPR100[10] , 
        \R_DATA_TEMPR101[10] , \R_DATA_TEMPR102[10] , 
        \R_DATA_TEMPR103[10] , \R_DATA_TEMPR104[10] , 
        \R_DATA_TEMPR105[10] , \R_DATA_TEMPR106[10] , 
        \R_DATA_TEMPR107[10] , \R_DATA_TEMPR108[10] , 
        \R_DATA_TEMPR109[10] , \R_DATA_TEMPR110[10] , 
        \R_DATA_TEMPR111[10] , \R_DATA_TEMPR112[10] , 
        \R_DATA_TEMPR113[10] , \R_DATA_TEMPR114[10] , 
        \R_DATA_TEMPR115[10] , \R_DATA_TEMPR116[10] , 
        \R_DATA_TEMPR117[10] , \R_DATA_TEMPR118[10] , 
        \R_DATA_TEMPR119[10] , \R_DATA_TEMPR120[10] , 
        \R_DATA_TEMPR121[10] , \R_DATA_TEMPR122[10] , 
        \R_DATA_TEMPR123[10] , \R_DATA_TEMPR124[10] , 
        \R_DATA_TEMPR125[10] , \R_DATA_TEMPR126[10] , 
        \R_DATA_TEMPR127[10] , \R_DATA_TEMPR0[11] , 
        \R_DATA_TEMPR1[11] , \R_DATA_TEMPR2[11] , \R_DATA_TEMPR3[11] , 
        \R_DATA_TEMPR4[11] , \R_DATA_TEMPR5[11] , \R_DATA_TEMPR6[11] , 
        \R_DATA_TEMPR7[11] , \R_DATA_TEMPR8[11] , \R_DATA_TEMPR9[11] , 
        \R_DATA_TEMPR10[11] , \R_DATA_TEMPR11[11] , 
        \R_DATA_TEMPR12[11] , \R_DATA_TEMPR13[11] , 
        \R_DATA_TEMPR14[11] , \R_DATA_TEMPR15[11] , 
        \R_DATA_TEMPR16[11] , \R_DATA_TEMPR17[11] , 
        \R_DATA_TEMPR18[11] , \R_DATA_TEMPR19[11] , 
        \R_DATA_TEMPR20[11] , \R_DATA_TEMPR21[11] , 
        \R_DATA_TEMPR22[11] , \R_DATA_TEMPR23[11] , 
        \R_DATA_TEMPR24[11] , \R_DATA_TEMPR25[11] , 
        \R_DATA_TEMPR26[11] , \R_DATA_TEMPR27[11] , 
        \R_DATA_TEMPR28[11] , \R_DATA_TEMPR29[11] , 
        \R_DATA_TEMPR30[11] , \R_DATA_TEMPR31[11] , 
        \R_DATA_TEMPR32[11] , \R_DATA_TEMPR33[11] , 
        \R_DATA_TEMPR34[11] , \R_DATA_TEMPR35[11] , 
        \R_DATA_TEMPR36[11] , \R_DATA_TEMPR37[11] , 
        \R_DATA_TEMPR38[11] , \R_DATA_TEMPR39[11] , 
        \R_DATA_TEMPR40[11] , \R_DATA_TEMPR41[11] , 
        \R_DATA_TEMPR42[11] , \R_DATA_TEMPR43[11] , 
        \R_DATA_TEMPR44[11] , \R_DATA_TEMPR45[11] , 
        \R_DATA_TEMPR46[11] , \R_DATA_TEMPR47[11] , 
        \R_DATA_TEMPR48[11] , \R_DATA_TEMPR49[11] , 
        \R_DATA_TEMPR50[11] , \R_DATA_TEMPR51[11] , 
        \R_DATA_TEMPR52[11] , \R_DATA_TEMPR53[11] , 
        \R_DATA_TEMPR54[11] , \R_DATA_TEMPR55[11] , 
        \R_DATA_TEMPR56[11] , \R_DATA_TEMPR57[11] , 
        \R_DATA_TEMPR58[11] , \R_DATA_TEMPR59[11] , 
        \R_DATA_TEMPR60[11] , \R_DATA_TEMPR61[11] , 
        \R_DATA_TEMPR62[11] , \R_DATA_TEMPR63[11] , 
        \R_DATA_TEMPR64[11] , \R_DATA_TEMPR65[11] , 
        \R_DATA_TEMPR66[11] , \R_DATA_TEMPR67[11] , 
        \R_DATA_TEMPR68[11] , \R_DATA_TEMPR69[11] , 
        \R_DATA_TEMPR70[11] , \R_DATA_TEMPR71[11] , 
        \R_DATA_TEMPR72[11] , \R_DATA_TEMPR73[11] , 
        \R_DATA_TEMPR74[11] , \R_DATA_TEMPR75[11] , 
        \R_DATA_TEMPR76[11] , \R_DATA_TEMPR77[11] , 
        \R_DATA_TEMPR78[11] , \R_DATA_TEMPR79[11] , 
        \R_DATA_TEMPR80[11] , \R_DATA_TEMPR81[11] , 
        \R_DATA_TEMPR82[11] , \R_DATA_TEMPR83[11] , 
        \R_DATA_TEMPR84[11] , \R_DATA_TEMPR85[11] , 
        \R_DATA_TEMPR86[11] , \R_DATA_TEMPR87[11] , 
        \R_DATA_TEMPR88[11] , \R_DATA_TEMPR89[11] , 
        \R_DATA_TEMPR90[11] , \R_DATA_TEMPR91[11] , 
        \R_DATA_TEMPR92[11] , \R_DATA_TEMPR93[11] , 
        \R_DATA_TEMPR94[11] , \R_DATA_TEMPR95[11] , 
        \R_DATA_TEMPR96[11] , \R_DATA_TEMPR97[11] , 
        \R_DATA_TEMPR98[11] , \R_DATA_TEMPR99[11] , 
        \R_DATA_TEMPR100[11] , \R_DATA_TEMPR101[11] , 
        \R_DATA_TEMPR102[11] , \R_DATA_TEMPR103[11] , 
        \R_DATA_TEMPR104[11] , \R_DATA_TEMPR105[11] , 
        \R_DATA_TEMPR106[11] , \R_DATA_TEMPR107[11] , 
        \R_DATA_TEMPR108[11] , \R_DATA_TEMPR109[11] , 
        \R_DATA_TEMPR110[11] , \R_DATA_TEMPR111[11] , 
        \R_DATA_TEMPR112[11] , \R_DATA_TEMPR113[11] , 
        \R_DATA_TEMPR114[11] , \R_DATA_TEMPR115[11] , 
        \R_DATA_TEMPR116[11] , \R_DATA_TEMPR117[11] , 
        \R_DATA_TEMPR118[11] , \R_DATA_TEMPR119[11] , 
        \R_DATA_TEMPR120[11] , \R_DATA_TEMPR121[11] , 
        \R_DATA_TEMPR122[11] , \R_DATA_TEMPR123[11] , 
        \R_DATA_TEMPR124[11] , \R_DATA_TEMPR125[11] , 
        \R_DATA_TEMPR126[11] , \R_DATA_TEMPR127[11] , 
        \R_DATA_TEMPR0[12] , \R_DATA_TEMPR1[12] , \R_DATA_TEMPR2[12] , 
        \R_DATA_TEMPR3[12] , \R_DATA_TEMPR4[12] , \R_DATA_TEMPR5[12] , 
        \R_DATA_TEMPR6[12] , \R_DATA_TEMPR7[12] , \R_DATA_TEMPR8[12] , 
        \R_DATA_TEMPR9[12] , \R_DATA_TEMPR10[12] , 
        \R_DATA_TEMPR11[12] , \R_DATA_TEMPR12[12] , 
        \R_DATA_TEMPR13[12] , \R_DATA_TEMPR14[12] , 
        \R_DATA_TEMPR15[12] , \R_DATA_TEMPR16[12] , 
        \R_DATA_TEMPR17[12] , \R_DATA_TEMPR18[12] , 
        \R_DATA_TEMPR19[12] , \R_DATA_TEMPR20[12] , 
        \R_DATA_TEMPR21[12] , \R_DATA_TEMPR22[12] , 
        \R_DATA_TEMPR23[12] , \R_DATA_TEMPR24[12] , 
        \R_DATA_TEMPR25[12] , \R_DATA_TEMPR26[12] , 
        \R_DATA_TEMPR27[12] , \R_DATA_TEMPR28[12] , 
        \R_DATA_TEMPR29[12] , \R_DATA_TEMPR30[12] , 
        \R_DATA_TEMPR31[12] , \R_DATA_TEMPR32[12] , 
        \R_DATA_TEMPR33[12] , \R_DATA_TEMPR34[12] , 
        \R_DATA_TEMPR35[12] , \R_DATA_TEMPR36[12] , 
        \R_DATA_TEMPR37[12] , \R_DATA_TEMPR38[12] , 
        \R_DATA_TEMPR39[12] , \R_DATA_TEMPR40[12] , 
        \R_DATA_TEMPR41[12] , \R_DATA_TEMPR42[12] , 
        \R_DATA_TEMPR43[12] , \R_DATA_TEMPR44[12] , 
        \R_DATA_TEMPR45[12] , \R_DATA_TEMPR46[12] , 
        \R_DATA_TEMPR47[12] , \R_DATA_TEMPR48[12] , 
        \R_DATA_TEMPR49[12] , \R_DATA_TEMPR50[12] , 
        \R_DATA_TEMPR51[12] , \R_DATA_TEMPR52[12] , 
        \R_DATA_TEMPR53[12] , \R_DATA_TEMPR54[12] , 
        \R_DATA_TEMPR55[12] , \R_DATA_TEMPR56[12] , 
        \R_DATA_TEMPR57[12] , \R_DATA_TEMPR58[12] , 
        \R_DATA_TEMPR59[12] , \R_DATA_TEMPR60[12] , 
        \R_DATA_TEMPR61[12] , \R_DATA_TEMPR62[12] , 
        \R_DATA_TEMPR63[12] , \R_DATA_TEMPR64[12] , 
        \R_DATA_TEMPR65[12] , \R_DATA_TEMPR66[12] , 
        \R_DATA_TEMPR67[12] , \R_DATA_TEMPR68[12] , 
        \R_DATA_TEMPR69[12] , \R_DATA_TEMPR70[12] , 
        \R_DATA_TEMPR71[12] , \R_DATA_TEMPR72[12] , 
        \R_DATA_TEMPR73[12] , \R_DATA_TEMPR74[12] , 
        \R_DATA_TEMPR75[12] , \R_DATA_TEMPR76[12] , 
        \R_DATA_TEMPR77[12] , \R_DATA_TEMPR78[12] , 
        \R_DATA_TEMPR79[12] , \R_DATA_TEMPR80[12] , 
        \R_DATA_TEMPR81[12] , \R_DATA_TEMPR82[12] , 
        \R_DATA_TEMPR83[12] , \R_DATA_TEMPR84[12] , 
        \R_DATA_TEMPR85[12] , \R_DATA_TEMPR86[12] , 
        \R_DATA_TEMPR87[12] , \R_DATA_TEMPR88[12] , 
        \R_DATA_TEMPR89[12] , \R_DATA_TEMPR90[12] , 
        \R_DATA_TEMPR91[12] , \R_DATA_TEMPR92[12] , 
        \R_DATA_TEMPR93[12] , \R_DATA_TEMPR94[12] , 
        \R_DATA_TEMPR95[12] , \R_DATA_TEMPR96[12] , 
        \R_DATA_TEMPR97[12] , \R_DATA_TEMPR98[12] , 
        \R_DATA_TEMPR99[12] , \R_DATA_TEMPR100[12] , 
        \R_DATA_TEMPR101[12] , \R_DATA_TEMPR102[12] , 
        \R_DATA_TEMPR103[12] , \R_DATA_TEMPR104[12] , 
        \R_DATA_TEMPR105[12] , \R_DATA_TEMPR106[12] , 
        \R_DATA_TEMPR107[12] , \R_DATA_TEMPR108[12] , 
        \R_DATA_TEMPR109[12] , \R_DATA_TEMPR110[12] , 
        \R_DATA_TEMPR111[12] , \R_DATA_TEMPR112[12] , 
        \R_DATA_TEMPR113[12] , \R_DATA_TEMPR114[12] , 
        \R_DATA_TEMPR115[12] , \R_DATA_TEMPR116[12] , 
        \R_DATA_TEMPR117[12] , \R_DATA_TEMPR118[12] , 
        \R_DATA_TEMPR119[12] , \R_DATA_TEMPR120[12] , 
        \R_DATA_TEMPR121[12] , \R_DATA_TEMPR122[12] , 
        \R_DATA_TEMPR123[12] , \R_DATA_TEMPR124[12] , 
        \R_DATA_TEMPR125[12] , \R_DATA_TEMPR126[12] , 
        \R_DATA_TEMPR127[12] , \R_DATA_TEMPR0[13] , 
        \R_DATA_TEMPR1[13] , \R_DATA_TEMPR2[13] , \R_DATA_TEMPR3[13] , 
        \R_DATA_TEMPR4[13] , \R_DATA_TEMPR5[13] , \R_DATA_TEMPR6[13] , 
        \R_DATA_TEMPR7[13] , \R_DATA_TEMPR8[13] , \R_DATA_TEMPR9[13] , 
        \R_DATA_TEMPR10[13] , \R_DATA_TEMPR11[13] , 
        \R_DATA_TEMPR12[13] , \R_DATA_TEMPR13[13] , 
        \R_DATA_TEMPR14[13] , \R_DATA_TEMPR15[13] , 
        \R_DATA_TEMPR16[13] , \R_DATA_TEMPR17[13] , 
        \R_DATA_TEMPR18[13] , \R_DATA_TEMPR19[13] , 
        \R_DATA_TEMPR20[13] , \R_DATA_TEMPR21[13] , 
        \R_DATA_TEMPR22[13] , \R_DATA_TEMPR23[13] , 
        \R_DATA_TEMPR24[13] , \R_DATA_TEMPR25[13] , 
        \R_DATA_TEMPR26[13] , \R_DATA_TEMPR27[13] , 
        \R_DATA_TEMPR28[13] , \R_DATA_TEMPR29[13] , 
        \R_DATA_TEMPR30[13] , \R_DATA_TEMPR31[13] , 
        \R_DATA_TEMPR32[13] , \R_DATA_TEMPR33[13] , 
        \R_DATA_TEMPR34[13] , \R_DATA_TEMPR35[13] , 
        \R_DATA_TEMPR36[13] , \R_DATA_TEMPR37[13] , 
        \R_DATA_TEMPR38[13] , \R_DATA_TEMPR39[13] , 
        \R_DATA_TEMPR40[13] , \R_DATA_TEMPR41[13] , 
        \R_DATA_TEMPR42[13] , \R_DATA_TEMPR43[13] , 
        \R_DATA_TEMPR44[13] , \R_DATA_TEMPR45[13] , 
        \R_DATA_TEMPR46[13] , \R_DATA_TEMPR47[13] , 
        \R_DATA_TEMPR48[13] , \R_DATA_TEMPR49[13] , 
        \R_DATA_TEMPR50[13] , \R_DATA_TEMPR51[13] , 
        \R_DATA_TEMPR52[13] , \R_DATA_TEMPR53[13] , 
        \R_DATA_TEMPR54[13] , \R_DATA_TEMPR55[13] , 
        \R_DATA_TEMPR56[13] , \R_DATA_TEMPR57[13] , 
        \R_DATA_TEMPR58[13] , \R_DATA_TEMPR59[13] , 
        \R_DATA_TEMPR60[13] , \R_DATA_TEMPR61[13] , 
        \R_DATA_TEMPR62[13] , \R_DATA_TEMPR63[13] , 
        \R_DATA_TEMPR64[13] , \R_DATA_TEMPR65[13] , 
        \R_DATA_TEMPR66[13] , \R_DATA_TEMPR67[13] , 
        \R_DATA_TEMPR68[13] , \R_DATA_TEMPR69[13] , 
        \R_DATA_TEMPR70[13] , \R_DATA_TEMPR71[13] , 
        \R_DATA_TEMPR72[13] , \R_DATA_TEMPR73[13] , 
        \R_DATA_TEMPR74[13] , \R_DATA_TEMPR75[13] , 
        \R_DATA_TEMPR76[13] , \R_DATA_TEMPR77[13] , 
        \R_DATA_TEMPR78[13] , \R_DATA_TEMPR79[13] , 
        \R_DATA_TEMPR80[13] , \R_DATA_TEMPR81[13] , 
        \R_DATA_TEMPR82[13] , \R_DATA_TEMPR83[13] , 
        \R_DATA_TEMPR84[13] , \R_DATA_TEMPR85[13] , 
        \R_DATA_TEMPR86[13] , \R_DATA_TEMPR87[13] , 
        \R_DATA_TEMPR88[13] , \R_DATA_TEMPR89[13] , 
        \R_DATA_TEMPR90[13] , \R_DATA_TEMPR91[13] , 
        \R_DATA_TEMPR92[13] , \R_DATA_TEMPR93[13] , 
        \R_DATA_TEMPR94[13] , \R_DATA_TEMPR95[13] , 
        \R_DATA_TEMPR96[13] , \R_DATA_TEMPR97[13] , 
        \R_DATA_TEMPR98[13] , \R_DATA_TEMPR99[13] , 
        \R_DATA_TEMPR100[13] , \R_DATA_TEMPR101[13] , 
        \R_DATA_TEMPR102[13] , \R_DATA_TEMPR103[13] , 
        \R_DATA_TEMPR104[13] , \R_DATA_TEMPR105[13] , 
        \R_DATA_TEMPR106[13] , \R_DATA_TEMPR107[13] , 
        \R_DATA_TEMPR108[13] , \R_DATA_TEMPR109[13] , 
        \R_DATA_TEMPR110[13] , \R_DATA_TEMPR111[13] , 
        \R_DATA_TEMPR112[13] , \R_DATA_TEMPR113[13] , 
        \R_DATA_TEMPR114[13] , \R_DATA_TEMPR115[13] , 
        \R_DATA_TEMPR116[13] , \R_DATA_TEMPR117[13] , 
        \R_DATA_TEMPR118[13] , \R_DATA_TEMPR119[13] , 
        \R_DATA_TEMPR120[13] , \R_DATA_TEMPR121[13] , 
        \R_DATA_TEMPR122[13] , \R_DATA_TEMPR123[13] , 
        \R_DATA_TEMPR124[13] , \R_DATA_TEMPR125[13] , 
        \R_DATA_TEMPR126[13] , \R_DATA_TEMPR127[13] , 
        \R_DATA_TEMPR0[14] , \R_DATA_TEMPR1[14] , \R_DATA_TEMPR2[14] , 
        \R_DATA_TEMPR3[14] , \R_DATA_TEMPR4[14] , \R_DATA_TEMPR5[14] , 
        \R_DATA_TEMPR6[14] , \R_DATA_TEMPR7[14] , \R_DATA_TEMPR8[14] , 
        \R_DATA_TEMPR9[14] , \R_DATA_TEMPR10[14] , 
        \R_DATA_TEMPR11[14] , \R_DATA_TEMPR12[14] , 
        \R_DATA_TEMPR13[14] , \R_DATA_TEMPR14[14] , 
        \R_DATA_TEMPR15[14] , \R_DATA_TEMPR16[14] , 
        \R_DATA_TEMPR17[14] , \R_DATA_TEMPR18[14] , 
        \R_DATA_TEMPR19[14] , \R_DATA_TEMPR20[14] , 
        \R_DATA_TEMPR21[14] , \R_DATA_TEMPR22[14] , 
        \R_DATA_TEMPR23[14] , \R_DATA_TEMPR24[14] , 
        \R_DATA_TEMPR25[14] , \R_DATA_TEMPR26[14] , 
        \R_DATA_TEMPR27[14] , \R_DATA_TEMPR28[14] , 
        \R_DATA_TEMPR29[14] , \R_DATA_TEMPR30[14] , 
        \R_DATA_TEMPR31[14] , \R_DATA_TEMPR32[14] , 
        \R_DATA_TEMPR33[14] , \R_DATA_TEMPR34[14] , 
        \R_DATA_TEMPR35[14] , \R_DATA_TEMPR36[14] , 
        \R_DATA_TEMPR37[14] , \R_DATA_TEMPR38[14] , 
        \R_DATA_TEMPR39[14] , \R_DATA_TEMPR40[14] , 
        \R_DATA_TEMPR41[14] , \R_DATA_TEMPR42[14] , 
        \R_DATA_TEMPR43[14] , \R_DATA_TEMPR44[14] , 
        \R_DATA_TEMPR45[14] , \R_DATA_TEMPR46[14] , 
        \R_DATA_TEMPR47[14] , \R_DATA_TEMPR48[14] , 
        \R_DATA_TEMPR49[14] , \R_DATA_TEMPR50[14] , 
        \R_DATA_TEMPR51[14] , \R_DATA_TEMPR52[14] , 
        \R_DATA_TEMPR53[14] , \R_DATA_TEMPR54[14] , 
        \R_DATA_TEMPR55[14] , \R_DATA_TEMPR56[14] , 
        \R_DATA_TEMPR57[14] , \R_DATA_TEMPR58[14] , 
        \R_DATA_TEMPR59[14] , \R_DATA_TEMPR60[14] , 
        \R_DATA_TEMPR61[14] , \R_DATA_TEMPR62[14] , 
        \R_DATA_TEMPR63[14] , \R_DATA_TEMPR64[14] , 
        \R_DATA_TEMPR65[14] , \R_DATA_TEMPR66[14] , 
        \R_DATA_TEMPR67[14] , \R_DATA_TEMPR68[14] , 
        \R_DATA_TEMPR69[14] , \R_DATA_TEMPR70[14] , 
        \R_DATA_TEMPR71[14] , \R_DATA_TEMPR72[14] , 
        \R_DATA_TEMPR73[14] , \R_DATA_TEMPR74[14] , 
        \R_DATA_TEMPR75[14] , \R_DATA_TEMPR76[14] , 
        \R_DATA_TEMPR77[14] , \R_DATA_TEMPR78[14] , 
        \R_DATA_TEMPR79[14] , \R_DATA_TEMPR80[14] , 
        \R_DATA_TEMPR81[14] , \R_DATA_TEMPR82[14] , 
        \R_DATA_TEMPR83[14] , \R_DATA_TEMPR84[14] , 
        \R_DATA_TEMPR85[14] , \R_DATA_TEMPR86[14] , 
        \R_DATA_TEMPR87[14] , \R_DATA_TEMPR88[14] , 
        \R_DATA_TEMPR89[14] , \R_DATA_TEMPR90[14] , 
        \R_DATA_TEMPR91[14] , \R_DATA_TEMPR92[14] , 
        \R_DATA_TEMPR93[14] , \R_DATA_TEMPR94[14] , 
        \R_DATA_TEMPR95[14] , \R_DATA_TEMPR96[14] , 
        \R_DATA_TEMPR97[14] , \R_DATA_TEMPR98[14] , 
        \R_DATA_TEMPR99[14] , \R_DATA_TEMPR100[14] , 
        \R_DATA_TEMPR101[14] , \R_DATA_TEMPR102[14] , 
        \R_DATA_TEMPR103[14] , \R_DATA_TEMPR104[14] , 
        \R_DATA_TEMPR105[14] , \R_DATA_TEMPR106[14] , 
        \R_DATA_TEMPR107[14] , \R_DATA_TEMPR108[14] , 
        \R_DATA_TEMPR109[14] , \R_DATA_TEMPR110[14] , 
        \R_DATA_TEMPR111[14] , \R_DATA_TEMPR112[14] , 
        \R_DATA_TEMPR113[14] , \R_DATA_TEMPR114[14] , 
        \R_DATA_TEMPR115[14] , \R_DATA_TEMPR116[14] , 
        \R_DATA_TEMPR117[14] , \R_DATA_TEMPR118[14] , 
        \R_DATA_TEMPR119[14] , \R_DATA_TEMPR120[14] , 
        \R_DATA_TEMPR121[14] , \R_DATA_TEMPR122[14] , 
        \R_DATA_TEMPR123[14] , \R_DATA_TEMPR124[14] , 
        \R_DATA_TEMPR125[14] , \R_DATA_TEMPR126[14] , 
        \R_DATA_TEMPR127[14] , \R_DATA_TEMPR0[15] , 
        \R_DATA_TEMPR1[15] , \R_DATA_TEMPR2[15] , \R_DATA_TEMPR3[15] , 
        \R_DATA_TEMPR4[15] , \R_DATA_TEMPR5[15] , \R_DATA_TEMPR6[15] , 
        \R_DATA_TEMPR7[15] , \R_DATA_TEMPR8[15] , \R_DATA_TEMPR9[15] , 
        \R_DATA_TEMPR10[15] , \R_DATA_TEMPR11[15] , 
        \R_DATA_TEMPR12[15] , \R_DATA_TEMPR13[15] , 
        \R_DATA_TEMPR14[15] , \R_DATA_TEMPR15[15] , 
        \R_DATA_TEMPR16[15] , \R_DATA_TEMPR17[15] , 
        \R_DATA_TEMPR18[15] , \R_DATA_TEMPR19[15] , 
        \R_DATA_TEMPR20[15] , \R_DATA_TEMPR21[15] , 
        \R_DATA_TEMPR22[15] , \R_DATA_TEMPR23[15] , 
        \R_DATA_TEMPR24[15] , \R_DATA_TEMPR25[15] , 
        \R_DATA_TEMPR26[15] , \R_DATA_TEMPR27[15] , 
        \R_DATA_TEMPR28[15] , \R_DATA_TEMPR29[15] , 
        \R_DATA_TEMPR30[15] , \R_DATA_TEMPR31[15] , 
        \R_DATA_TEMPR32[15] , \R_DATA_TEMPR33[15] , 
        \R_DATA_TEMPR34[15] , \R_DATA_TEMPR35[15] , 
        \R_DATA_TEMPR36[15] , \R_DATA_TEMPR37[15] , 
        \R_DATA_TEMPR38[15] , \R_DATA_TEMPR39[15] , 
        \R_DATA_TEMPR40[15] , \R_DATA_TEMPR41[15] , 
        \R_DATA_TEMPR42[15] , \R_DATA_TEMPR43[15] , 
        \R_DATA_TEMPR44[15] , \R_DATA_TEMPR45[15] , 
        \R_DATA_TEMPR46[15] , \R_DATA_TEMPR47[15] , 
        \R_DATA_TEMPR48[15] , \R_DATA_TEMPR49[15] , 
        \R_DATA_TEMPR50[15] , \R_DATA_TEMPR51[15] , 
        \R_DATA_TEMPR52[15] , \R_DATA_TEMPR53[15] , 
        \R_DATA_TEMPR54[15] , \R_DATA_TEMPR55[15] , 
        \R_DATA_TEMPR56[15] , \R_DATA_TEMPR57[15] , 
        \R_DATA_TEMPR58[15] , \R_DATA_TEMPR59[15] , 
        \R_DATA_TEMPR60[15] , \R_DATA_TEMPR61[15] , 
        \R_DATA_TEMPR62[15] , \R_DATA_TEMPR63[15] , 
        \R_DATA_TEMPR64[15] , \R_DATA_TEMPR65[15] , 
        \R_DATA_TEMPR66[15] , \R_DATA_TEMPR67[15] , 
        \R_DATA_TEMPR68[15] , \R_DATA_TEMPR69[15] , 
        \R_DATA_TEMPR70[15] , \R_DATA_TEMPR71[15] , 
        \R_DATA_TEMPR72[15] , \R_DATA_TEMPR73[15] , 
        \R_DATA_TEMPR74[15] , \R_DATA_TEMPR75[15] , 
        \R_DATA_TEMPR76[15] , \R_DATA_TEMPR77[15] , 
        \R_DATA_TEMPR78[15] , \R_DATA_TEMPR79[15] , 
        \R_DATA_TEMPR80[15] , \R_DATA_TEMPR81[15] , 
        \R_DATA_TEMPR82[15] , \R_DATA_TEMPR83[15] , 
        \R_DATA_TEMPR84[15] , \R_DATA_TEMPR85[15] , 
        \R_DATA_TEMPR86[15] , \R_DATA_TEMPR87[15] , 
        \R_DATA_TEMPR88[15] , \R_DATA_TEMPR89[15] , 
        \R_DATA_TEMPR90[15] , \R_DATA_TEMPR91[15] , 
        \R_DATA_TEMPR92[15] , \R_DATA_TEMPR93[15] , 
        \R_DATA_TEMPR94[15] , \R_DATA_TEMPR95[15] , 
        \R_DATA_TEMPR96[15] , \R_DATA_TEMPR97[15] , 
        \R_DATA_TEMPR98[15] , \R_DATA_TEMPR99[15] , 
        \R_DATA_TEMPR100[15] , \R_DATA_TEMPR101[15] , 
        \R_DATA_TEMPR102[15] , \R_DATA_TEMPR103[15] , 
        \R_DATA_TEMPR104[15] , \R_DATA_TEMPR105[15] , 
        \R_DATA_TEMPR106[15] , \R_DATA_TEMPR107[15] , 
        \R_DATA_TEMPR108[15] , \R_DATA_TEMPR109[15] , 
        \R_DATA_TEMPR110[15] , \R_DATA_TEMPR111[15] , 
        \R_DATA_TEMPR112[15] , \R_DATA_TEMPR113[15] , 
        \R_DATA_TEMPR114[15] , \R_DATA_TEMPR115[15] , 
        \R_DATA_TEMPR116[15] , \R_DATA_TEMPR117[15] , 
        \R_DATA_TEMPR118[15] , \R_DATA_TEMPR119[15] , 
        \R_DATA_TEMPR120[15] , \R_DATA_TEMPR121[15] , 
        \R_DATA_TEMPR122[15] , \R_DATA_TEMPR123[15] , 
        \R_DATA_TEMPR124[15] , \R_DATA_TEMPR125[15] , 
        \R_DATA_TEMPR126[15] , \R_DATA_TEMPR127[15] , 
        \R_DATA_TEMPR0[16] , \R_DATA_TEMPR1[16] , \R_DATA_TEMPR2[16] , 
        \R_DATA_TEMPR3[16] , \R_DATA_TEMPR4[16] , \R_DATA_TEMPR5[16] , 
        \R_DATA_TEMPR6[16] , \R_DATA_TEMPR7[16] , \R_DATA_TEMPR8[16] , 
        \R_DATA_TEMPR9[16] , \R_DATA_TEMPR10[16] , 
        \R_DATA_TEMPR11[16] , \R_DATA_TEMPR12[16] , 
        \R_DATA_TEMPR13[16] , \R_DATA_TEMPR14[16] , 
        \R_DATA_TEMPR15[16] , \R_DATA_TEMPR16[16] , 
        \R_DATA_TEMPR17[16] , \R_DATA_TEMPR18[16] , 
        \R_DATA_TEMPR19[16] , \R_DATA_TEMPR20[16] , 
        \R_DATA_TEMPR21[16] , \R_DATA_TEMPR22[16] , 
        \R_DATA_TEMPR23[16] , \R_DATA_TEMPR24[16] , 
        \R_DATA_TEMPR25[16] , \R_DATA_TEMPR26[16] , 
        \R_DATA_TEMPR27[16] , \R_DATA_TEMPR28[16] , 
        \R_DATA_TEMPR29[16] , \R_DATA_TEMPR30[16] , 
        \R_DATA_TEMPR31[16] , \R_DATA_TEMPR32[16] , 
        \R_DATA_TEMPR33[16] , \R_DATA_TEMPR34[16] , 
        \R_DATA_TEMPR35[16] , \R_DATA_TEMPR36[16] , 
        \R_DATA_TEMPR37[16] , \R_DATA_TEMPR38[16] , 
        \R_DATA_TEMPR39[16] , \R_DATA_TEMPR40[16] , 
        \R_DATA_TEMPR41[16] , \R_DATA_TEMPR42[16] , 
        \R_DATA_TEMPR43[16] , \R_DATA_TEMPR44[16] , 
        \R_DATA_TEMPR45[16] , \R_DATA_TEMPR46[16] , 
        \R_DATA_TEMPR47[16] , \R_DATA_TEMPR48[16] , 
        \R_DATA_TEMPR49[16] , \R_DATA_TEMPR50[16] , 
        \R_DATA_TEMPR51[16] , \R_DATA_TEMPR52[16] , 
        \R_DATA_TEMPR53[16] , \R_DATA_TEMPR54[16] , 
        \R_DATA_TEMPR55[16] , \R_DATA_TEMPR56[16] , 
        \R_DATA_TEMPR57[16] , \R_DATA_TEMPR58[16] , 
        \R_DATA_TEMPR59[16] , \R_DATA_TEMPR60[16] , 
        \R_DATA_TEMPR61[16] , \R_DATA_TEMPR62[16] , 
        \R_DATA_TEMPR63[16] , \R_DATA_TEMPR64[16] , 
        \R_DATA_TEMPR65[16] , \R_DATA_TEMPR66[16] , 
        \R_DATA_TEMPR67[16] , \R_DATA_TEMPR68[16] , 
        \R_DATA_TEMPR69[16] , \R_DATA_TEMPR70[16] , 
        \R_DATA_TEMPR71[16] , \R_DATA_TEMPR72[16] , 
        \R_DATA_TEMPR73[16] , \R_DATA_TEMPR74[16] , 
        \R_DATA_TEMPR75[16] , \R_DATA_TEMPR76[16] , 
        \R_DATA_TEMPR77[16] , \R_DATA_TEMPR78[16] , 
        \R_DATA_TEMPR79[16] , \R_DATA_TEMPR80[16] , 
        \R_DATA_TEMPR81[16] , \R_DATA_TEMPR82[16] , 
        \R_DATA_TEMPR83[16] , \R_DATA_TEMPR84[16] , 
        \R_DATA_TEMPR85[16] , \R_DATA_TEMPR86[16] , 
        \R_DATA_TEMPR87[16] , \R_DATA_TEMPR88[16] , 
        \R_DATA_TEMPR89[16] , \R_DATA_TEMPR90[16] , 
        \R_DATA_TEMPR91[16] , \R_DATA_TEMPR92[16] , 
        \R_DATA_TEMPR93[16] , \R_DATA_TEMPR94[16] , 
        \R_DATA_TEMPR95[16] , \R_DATA_TEMPR96[16] , 
        \R_DATA_TEMPR97[16] , \R_DATA_TEMPR98[16] , 
        \R_DATA_TEMPR99[16] , \R_DATA_TEMPR100[16] , 
        \R_DATA_TEMPR101[16] , \R_DATA_TEMPR102[16] , 
        \R_DATA_TEMPR103[16] , \R_DATA_TEMPR104[16] , 
        \R_DATA_TEMPR105[16] , \R_DATA_TEMPR106[16] , 
        \R_DATA_TEMPR107[16] , \R_DATA_TEMPR108[16] , 
        \R_DATA_TEMPR109[16] , \R_DATA_TEMPR110[16] , 
        \R_DATA_TEMPR111[16] , \R_DATA_TEMPR112[16] , 
        \R_DATA_TEMPR113[16] , \R_DATA_TEMPR114[16] , 
        \R_DATA_TEMPR115[16] , \R_DATA_TEMPR116[16] , 
        \R_DATA_TEMPR117[16] , \R_DATA_TEMPR118[16] , 
        \R_DATA_TEMPR119[16] , \R_DATA_TEMPR120[16] , 
        \R_DATA_TEMPR121[16] , \R_DATA_TEMPR122[16] , 
        \R_DATA_TEMPR123[16] , \R_DATA_TEMPR124[16] , 
        \R_DATA_TEMPR125[16] , \R_DATA_TEMPR126[16] , 
        \R_DATA_TEMPR127[16] , \R_DATA_TEMPR0[17] , 
        \R_DATA_TEMPR1[17] , \R_DATA_TEMPR2[17] , \R_DATA_TEMPR3[17] , 
        \R_DATA_TEMPR4[17] , \R_DATA_TEMPR5[17] , \R_DATA_TEMPR6[17] , 
        \R_DATA_TEMPR7[17] , \R_DATA_TEMPR8[17] , \R_DATA_TEMPR9[17] , 
        \R_DATA_TEMPR10[17] , \R_DATA_TEMPR11[17] , 
        \R_DATA_TEMPR12[17] , \R_DATA_TEMPR13[17] , 
        \R_DATA_TEMPR14[17] , \R_DATA_TEMPR15[17] , 
        \R_DATA_TEMPR16[17] , \R_DATA_TEMPR17[17] , 
        \R_DATA_TEMPR18[17] , \R_DATA_TEMPR19[17] , 
        \R_DATA_TEMPR20[17] , \R_DATA_TEMPR21[17] , 
        \R_DATA_TEMPR22[17] , \R_DATA_TEMPR23[17] , 
        \R_DATA_TEMPR24[17] , \R_DATA_TEMPR25[17] , 
        \R_DATA_TEMPR26[17] , \R_DATA_TEMPR27[17] , 
        \R_DATA_TEMPR28[17] , \R_DATA_TEMPR29[17] , 
        \R_DATA_TEMPR30[17] , \R_DATA_TEMPR31[17] , 
        \R_DATA_TEMPR32[17] , \R_DATA_TEMPR33[17] , 
        \R_DATA_TEMPR34[17] , \R_DATA_TEMPR35[17] , 
        \R_DATA_TEMPR36[17] , \R_DATA_TEMPR37[17] , 
        \R_DATA_TEMPR38[17] , \R_DATA_TEMPR39[17] , 
        \R_DATA_TEMPR40[17] , \R_DATA_TEMPR41[17] , 
        \R_DATA_TEMPR42[17] , \R_DATA_TEMPR43[17] , 
        \R_DATA_TEMPR44[17] , \R_DATA_TEMPR45[17] , 
        \R_DATA_TEMPR46[17] , \R_DATA_TEMPR47[17] , 
        \R_DATA_TEMPR48[17] , \R_DATA_TEMPR49[17] , 
        \R_DATA_TEMPR50[17] , \R_DATA_TEMPR51[17] , 
        \R_DATA_TEMPR52[17] , \R_DATA_TEMPR53[17] , 
        \R_DATA_TEMPR54[17] , \R_DATA_TEMPR55[17] , 
        \R_DATA_TEMPR56[17] , \R_DATA_TEMPR57[17] , 
        \R_DATA_TEMPR58[17] , \R_DATA_TEMPR59[17] , 
        \R_DATA_TEMPR60[17] , \R_DATA_TEMPR61[17] , 
        \R_DATA_TEMPR62[17] , \R_DATA_TEMPR63[17] , 
        \R_DATA_TEMPR64[17] , \R_DATA_TEMPR65[17] , 
        \R_DATA_TEMPR66[17] , \R_DATA_TEMPR67[17] , 
        \R_DATA_TEMPR68[17] , \R_DATA_TEMPR69[17] , 
        \R_DATA_TEMPR70[17] , \R_DATA_TEMPR71[17] , 
        \R_DATA_TEMPR72[17] , \R_DATA_TEMPR73[17] , 
        \R_DATA_TEMPR74[17] , \R_DATA_TEMPR75[17] , 
        \R_DATA_TEMPR76[17] , \R_DATA_TEMPR77[17] , 
        \R_DATA_TEMPR78[17] , \R_DATA_TEMPR79[17] , 
        \R_DATA_TEMPR80[17] , \R_DATA_TEMPR81[17] , 
        \R_DATA_TEMPR82[17] , \R_DATA_TEMPR83[17] , 
        \R_DATA_TEMPR84[17] , \R_DATA_TEMPR85[17] , 
        \R_DATA_TEMPR86[17] , \R_DATA_TEMPR87[17] , 
        \R_DATA_TEMPR88[17] , \R_DATA_TEMPR89[17] , 
        \R_DATA_TEMPR90[17] , \R_DATA_TEMPR91[17] , 
        \R_DATA_TEMPR92[17] , \R_DATA_TEMPR93[17] , 
        \R_DATA_TEMPR94[17] , \R_DATA_TEMPR95[17] , 
        \R_DATA_TEMPR96[17] , \R_DATA_TEMPR97[17] , 
        \R_DATA_TEMPR98[17] , \R_DATA_TEMPR99[17] , 
        \R_DATA_TEMPR100[17] , \R_DATA_TEMPR101[17] , 
        \R_DATA_TEMPR102[17] , \R_DATA_TEMPR103[17] , 
        \R_DATA_TEMPR104[17] , \R_DATA_TEMPR105[17] , 
        \R_DATA_TEMPR106[17] , \R_DATA_TEMPR107[17] , 
        \R_DATA_TEMPR108[17] , \R_DATA_TEMPR109[17] , 
        \R_DATA_TEMPR110[17] , \R_DATA_TEMPR111[17] , 
        \R_DATA_TEMPR112[17] , \R_DATA_TEMPR113[17] , 
        \R_DATA_TEMPR114[17] , \R_DATA_TEMPR115[17] , 
        \R_DATA_TEMPR116[17] , \R_DATA_TEMPR117[17] , 
        \R_DATA_TEMPR118[17] , \R_DATA_TEMPR119[17] , 
        \R_DATA_TEMPR120[17] , \R_DATA_TEMPR121[17] , 
        \R_DATA_TEMPR122[17] , \R_DATA_TEMPR123[17] , 
        \R_DATA_TEMPR124[17] , \R_DATA_TEMPR125[17] , 
        \R_DATA_TEMPR126[17] , \R_DATA_TEMPR127[17] , 
        \R_DATA_TEMPR0[18] , \R_DATA_TEMPR1[18] , \R_DATA_TEMPR2[18] , 
        \R_DATA_TEMPR3[18] , \R_DATA_TEMPR4[18] , \R_DATA_TEMPR5[18] , 
        \R_DATA_TEMPR6[18] , \R_DATA_TEMPR7[18] , \R_DATA_TEMPR8[18] , 
        \R_DATA_TEMPR9[18] , \R_DATA_TEMPR10[18] , 
        \R_DATA_TEMPR11[18] , \R_DATA_TEMPR12[18] , 
        \R_DATA_TEMPR13[18] , \R_DATA_TEMPR14[18] , 
        \R_DATA_TEMPR15[18] , \R_DATA_TEMPR16[18] , 
        \R_DATA_TEMPR17[18] , \R_DATA_TEMPR18[18] , 
        \R_DATA_TEMPR19[18] , \R_DATA_TEMPR20[18] , 
        \R_DATA_TEMPR21[18] , \R_DATA_TEMPR22[18] , 
        \R_DATA_TEMPR23[18] , \R_DATA_TEMPR24[18] , 
        \R_DATA_TEMPR25[18] , \R_DATA_TEMPR26[18] , 
        \R_DATA_TEMPR27[18] , \R_DATA_TEMPR28[18] , 
        \R_DATA_TEMPR29[18] , \R_DATA_TEMPR30[18] , 
        \R_DATA_TEMPR31[18] , \R_DATA_TEMPR32[18] , 
        \R_DATA_TEMPR33[18] , \R_DATA_TEMPR34[18] , 
        \R_DATA_TEMPR35[18] , \R_DATA_TEMPR36[18] , 
        \R_DATA_TEMPR37[18] , \R_DATA_TEMPR38[18] , 
        \R_DATA_TEMPR39[18] , \R_DATA_TEMPR40[18] , 
        \R_DATA_TEMPR41[18] , \R_DATA_TEMPR42[18] , 
        \R_DATA_TEMPR43[18] , \R_DATA_TEMPR44[18] , 
        \R_DATA_TEMPR45[18] , \R_DATA_TEMPR46[18] , 
        \R_DATA_TEMPR47[18] , \R_DATA_TEMPR48[18] , 
        \R_DATA_TEMPR49[18] , \R_DATA_TEMPR50[18] , 
        \R_DATA_TEMPR51[18] , \R_DATA_TEMPR52[18] , 
        \R_DATA_TEMPR53[18] , \R_DATA_TEMPR54[18] , 
        \R_DATA_TEMPR55[18] , \R_DATA_TEMPR56[18] , 
        \R_DATA_TEMPR57[18] , \R_DATA_TEMPR58[18] , 
        \R_DATA_TEMPR59[18] , \R_DATA_TEMPR60[18] , 
        \R_DATA_TEMPR61[18] , \R_DATA_TEMPR62[18] , 
        \R_DATA_TEMPR63[18] , \R_DATA_TEMPR64[18] , 
        \R_DATA_TEMPR65[18] , \R_DATA_TEMPR66[18] , 
        \R_DATA_TEMPR67[18] , \R_DATA_TEMPR68[18] , 
        \R_DATA_TEMPR69[18] , \R_DATA_TEMPR70[18] , 
        \R_DATA_TEMPR71[18] , \R_DATA_TEMPR72[18] , 
        \R_DATA_TEMPR73[18] , \R_DATA_TEMPR74[18] , 
        \R_DATA_TEMPR75[18] , \R_DATA_TEMPR76[18] , 
        \R_DATA_TEMPR77[18] , \R_DATA_TEMPR78[18] , 
        \R_DATA_TEMPR79[18] , \R_DATA_TEMPR80[18] , 
        \R_DATA_TEMPR81[18] , \R_DATA_TEMPR82[18] , 
        \R_DATA_TEMPR83[18] , \R_DATA_TEMPR84[18] , 
        \R_DATA_TEMPR85[18] , \R_DATA_TEMPR86[18] , 
        \R_DATA_TEMPR87[18] , \R_DATA_TEMPR88[18] , 
        \R_DATA_TEMPR89[18] , \R_DATA_TEMPR90[18] , 
        \R_DATA_TEMPR91[18] , \R_DATA_TEMPR92[18] , 
        \R_DATA_TEMPR93[18] , \R_DATA_TEMPR94[18] , 
        \R_DATA_TEMPR95[18] , \R_DATA_TEMPR96[18] , 
        \R_DATA_TEMPR97[18] , \R_DATA_TEMPR98[18] , 
        \R_DATA_TEMPR99[18] , \R_DATA_TEMPR100[18] , 
        \R_DATA_TEMPR101[18] , \R_DATA_TEMPR102[18] , 
        \R_DATA_TEMPR103[18] , \R_DATA_TEMPR104[18] , 
        \R_DATA_TEMPR105[18] , \R_DATA_TEMPR106[18] , 
        \R_DATA_TEMPR107[18] , \R_DATA_TEMPR108[18] , 
        \R_DATA_TEMPR109[18] , \R_DATA_TEMPR110[18] , 
        \R_DATA_TEMPR111[18] , \R_DATA_TEMPR112[18] , 
        \R_DATA_TEMPR113[18] , \R_DATA_TEMPR114[18] , 
        \R_DATA_TEMPR115[18] , \R_DATA_TEMPR116[18] , 
        \R_DATA_TEMPR117[18] , \R_DATA_TEMPR118[18] , 
        \R_DATA_TEMPR119[18] , \R_DATA_TEMPR120[18] , 
        \R_DATA_TEMPR121[18] , \R_DATA_TEMPR122[18] , 
        \R_DATA_TEMPR123[18] , \R_DATA_TEMPR124[18] , 
        \R_DATA_TEMPR125[18] , \R_DATA_TEMPR126[18] , 
        \R_DATA_TEMPR127[18] , \R_DATA_TEMPR0[19] , 
        \R_DATA_TEMPR1[19] , \R_DATA_TEMPR2[19] , \R_DATA_TEMPR3[19] , 
        \R_DATA_TEMPR4[19] , \R_DATA_TEMPR5[19] , \R_DATA_TEMPR6[19] , 
        \R_DATA_TEMPR7[19] , \R_DATA_TEMPR8[19] , \R_DATA_TEMPR9[19] , 
        \R_DATA_TEMPR10[19] , \R_DATA_TEMPR11[19] , 
        \R_DATA_TEMPR12[19] , \R_DATA_TEMPR13[19] , 
        \R_DATA_TEMPR14[19] , \R_DATA_TEMPR15[19] , 
        \R_DATA_TEMPR16[19] , \R_DATA_TEMPR17[19] , 
        \R_DATA_TEMPR18[19] , \R_DATA_TEMPR19[19] , 
        \R_DATA_TEMPR20[19] , \R_DATA_TEMPR21[19] , 
        \R_DATA_TEMPR22[19] , \R_DATA_TEMPR23[19] , 
        \R_DATA_TEMPR24[19] , \R_DATA_TEMPR25[19] , 
        \R_DATA_TEMPR26[19] , \R_DATA_TEMPR27[19] , 
        \R_DATA_TEMPR28[19] , \R_DATA_TEMPR29[19] , 
        \R_DATA_TEMPR30[19] , \R_DATA_TEMPR31[19] , 
        \R_DATA_TEMPR32[19] , \R_DATA_TEMPR33[19] , 
        \R_DATA_TEMPR34[19] , \R_DATA_TEMPR35[19] , 
        \R_DATA_TEMPR36[19] , \R_DATA_TEMPR37[19] , 
        \R_DATA_TEMPR38[19] , \R_DATA_TEMPR39[19] , 
        \R_DATA_TEMPR40[19] , \R_DATA_TEMPR41[19] , 
        \R_DATA_TEMPR42[19] , \R_DATA_TEMPR43[19] , 
        \R_DATA_TEMPR44[19] , \R_DATA_TEMPR45[19] , 
        \R_DATA_TEMPR46[19] , \R_DATA_TEMPR47[19] , 
        \R_DATA_TEMPR48[19] , \R_DATA_TEMPR49[19] , 
        \R_DATA_TEMPR50[19] , \R_DATA_TEMPR51[19] , 
        \R_DATA_TEMPR52[19] , \R_DATA_TEMPR53[19] , 
        \R_DATA_TEMPR54[19] , \R_DATA_TEMPR55[19] , 
        \R_DATA_TEMPR56[19] , \R_DATA_TEMPR57[19] , 
        \R_DATA_TEMPR58[19] , \R_DATA_TEMPR59[19] , 
        \R_DATA_TEMPR60[19] , \R_DATA_TEMPR61[19] , 
        \R_DATA_TEMPR62[19] , \R_DATA_TEMPR63[19] , 
        \R_DATA_TEMPR64[19] , \R_DATA_TEMPR65[19] , 
        \R_DATA_TEMPR66[19] , \R_DATA_TEMPR67[19] , 
        \R_DATA_TEMPR68[19] , \R_DATA_TEMPR69[19] , 
        \R_DATA_TEMPR70[19] , \R_DATA_TEMPR71[19] , 
        \R_DATA_TEMPR72[19] , \R_DATA_TEMPR73[19] , 
        \R_DATA_TEMPR74[19] , \R_DATA_TEMPR75[19] , 
        \R_DATA_TEMPR76[19] , \R_DATA_TEMPR77[19] , 
        \R_DATA_TEMPR78[19] , \R_DATA_TEMPR79[19] , 
        \R_DATA_TEMPR80[19] , \R_DATA_TEMPR81[19] , 
        \R_DATA_TEMPR82[19] , \R_DATA_TEMPR83[19] , 
        \R_DATA_TEMPR84[19] , \R_DATA_TEMPR85[19] , 
        \R_DATA_TEMPR86[19] , \R_DATA_TEMPR87[19] , 
        \R_DATA_TEMPR88[19] , \R_DATA_TEMPR89[19] , 
        \R_DATA_TEMPR90[19] , \R_DATA_TEMPR91[19] , 
        \R_DATA_TEMPR92[19] , \R_DATA_TEMPR93[19] , 
        \R_DATA_TEMPR94[19] , \R_DATA_TEMPR95[19] , 
        \R_DATA_TEMPR96[19] , \R_DATA_TEMPR97[19] , 
        \R_DATA_TEMPR98[19] , \R_DATA_TEMPR99[19] , 
        \R_DATA_TEMPR100[19] , \R_DATA_TEMPR101[19] , 
        \R_DATA_TEMPR102[19] , \R_DATA_TEMPR103[19] , 
        \R_DATA_TEMPR104[19] , \R_DATA_TEMPR105[19] , 
        \R_DATA_TEMPR106[19] , \R_DATA_TEMPR107[19] , 
        \R_DATA_TEMPR108[19] , \R_DATA_TEMPR109[19] , 
        \R_DATA_TEMPR110[19] , \R_DATA_TEMPR111[19] , 
        \R_DATA_TEMPR112[19] , \R_DATA_TEMPR113[19] , 
        \R_DATA_TEMPR114[19] , \R_DATA_TEMPR115[19] , 
        \R_DATA_TEMPR116[19] , \R_DATA_TEMPR117[19] , 
        \R_DATA_TEMPR118[19] , \R_DATA_TEMPR119[19] , 
        \R_DATA_TEMPR120[19] , \R_DATA_TEMPR121[19] , 
        \R_DATA_TEMPR122[19] , \R_DATA_TEMPR123[19] , 
        \R_DATA_TEMPR124[19] , \R_DATA_TEMPR125[19] , 
        \R_DATA_TEMPR126[19] , \R_DATA_TEMPR127[19] , 
        \R_DATA_TEMPR0[20] , \R_DATA_TEMPR1[20] , \R_DATA_TEMPR2[20] , 
        \R_DATA_TEMPR3[20] , \R_DATA_TEMPR4[20] , \R_DATA_TEMPR5[20] , 
        \R_DATA_TEMPR6[20] , \R_DATA_TEMPR7[20] , \R_DATA_TEMPR8[20] , 
        \R_DATA_TEMPR9[20] , \R_DATA_TEMPR10[20] , 
        \R_DATA_TEMPR11[20] , \R_DATA_TEMPR12[20] , 
        \R_DATA_TEMPR13[20] , \R_DATA_TEMPR14[20] , 
        \R_DATA_TEMPR15[20] , \R_DATA_TEMPR16[20] , 
        \R_DATA_TEMPR17[20] , \R_DATA_TEMPR18[20] , 
        \R_DATA_TEMPR19[20] , \R_DATA_TEMPR20[20] , 
        \R_DATA_TEMPR21[20] , \R_DATA_TEMPR22[20] , 
        \R_DATA_TEMPR23[20] , \R_DATA_TEMPR24[20] , 
        \R_DATA_TEMPR25[20] , \R_DATA_TEMPR26[20] , 
        \R_DATA_TEMPR27[20] , \R_DATA_TEMPR28[20] , 
        \R_DATA_TEMPR29[20] , \R_DATA_TEMPR30[20] , 
        \R_DATA_TEMPR31[20] , \R_DATA_TEMPR32[20] , 
        \R_DATA_TEMPR33[20] , \R_DATA_TEMPR34[20] , 
        \R_DATA_TEMPR35[20] , \R_DATA_TEMPR36[20] , 
        \R_DATA_TEMPR37[20] , \R_DATA_TEMPR38[20] , 
        \R_DATA_TEMPR39[20] , \R_DATA_TEMPR40[20] , 
        \R_DATA_TEMPR41[20] , \R_DATA_TEMPR42[20] , 
        \R_DATA_TEMPR43[20] , \R_DATA_TEMPR44[20] , 
        \R_DATA_TEMPR45[20] , \R_DATA_TEMPR46[20] , 
        \R_DATA_TEMPR47[20] , \R_DATA_TEMPR48[20] , 
        \R_DATA_TEMPR49[20] , \R_DATA_TEMPR50[20] , 
        \R_DATA_TEMPR51[20] , \R_DATA_TEMPR52[20] , 
        \R_DATA_TEMPR53[20] , \R_DATA_TEMPR54[20] , 
        \R_DATA_TEMPR55[20] , \R_DATA_TEMPR56[20] , 
        \R_DATA_TEMPR57[20] , \R_DATA_TEMPR58[20] , 
        \R_DATA_TEMPR59[20] , \R_DATA_TEMPR60[20] , 
        \R_DATA_TEMPR61[20] , \R_DATA_TEMPR62[20] , 
        \R_DATA_TEMPR63[20] , \R_DATA_TEMPR64[20] , 
        \R_DATA_TEMPR65[20] , \R_DATA_TEMPR66[20] , 
        \R_DATA_TEMPR67[20] , \R_DATA_TEMPR68[20] , 
        \R_DATA_TEMPR69[20] , \R_DATA_TEMPR70[20] , 
        \R_DATA_TEMPR71[20] , \R_DATA_TEMPR72[20] , 
        \R_DATA_TEMPR73[20] , \R_DATA_TEMPR74[20] , 
        \R_DATA_TEMPR75[20] , \R_DATA_TEMPR76[20] , 
        \R_DATA_TEMPR77[20] , \R_DATA_TEMPR78[20] , 
        \R_DATA_TEMPR79[20] , \R_DATA_TEMPR80[20] , 
        \R_DATA_TEMPR81[20] , \R_DATA_TEMPR82[20] , 
        \R_DATA_TEMPR83[20] , \R_DATA_TEMPR84[20] , 
        \R_DATA_TEMPR85[20] , \R_DATA_TEMPR86[20] , 
        \R_DATA_TEMPR87[20] , \R_DATA_TEMPR88[20] , 
        \R_DATA_TEMPR89[20] , \R_DATA_TEMPR90[20] , 
        \R_DATA_TEMPR91[20] , \R_DATA_TEMPR92[20] , 
        \R_DATA_TEMPR93[20] , \R_DATA_TEMPR94[20] , 
        \R_DATA_TEMPR95[20] , \R_DATA_TEMPR96[20] , 
        \R_DATA_TEMPR97[20] , \R_DATA_TEMPR98[20] , 
        \R_DATA_TEMPR99[20] , \R_DATA_TEMPR100[20] , 
        \R_DATA_TEMPR101[20] , \R_DATA_TEMPR102[20] , 
        \R_DATA_TEMPR103[20] , \R_DATA_TEMPR104[20] , 
        \R_DATA_TEMPR105[20] , \R_DATA_TEMPR106[20] , 
        \R_DATA_TEMPR107[20] , \R_DATA_TEMPR108[20] , 
        \R_DATA_TEMPR109[20] , \R_DATA_TEMPR110[20] , 
        \R_DATA_TEMPR111[20] , \R_DATA_TEMPR112[20] , 
        \R_DATA_TEMPR113[20] , \R_DATA_TEMPR114[20] , 
        \R_DATA_TEMPR115[20] , \R_DATA_TEMPR116[20] , 
        \R_DATA_TEMPR117[20] , \R_DATA_TEMPR118[20] , 
        \R_DATA_TEMPR119[20] , \R_DATA_TEMPR120[20] , 
        \R_DATA_TEMPR121[20] , \R_DATA_TEMPR122[20] , 
        \R_DATA_TEMPR123[20] , \R_DATA_TEMPR124[20] , 
        \R_DATA_TEMPR125[20] , \R_DATA_TEMPR126[20] , 
        \R_DATA_TEMPR127[20] , \R_DATA_TEMPR0[21] , 
        \R_DATA_TEMPR1[21] , \R_DATA_TEMPR2[21] , \R_DATA_TEMPR3[21] , 
        \R_DATA_TEMPR4[21] , \R_DATA_TEMPR5[21] , \R_DATA_TEMPR6[21] , 
        \R_DATA_TEMPR7[21] , \R_DATA_TEMPR8[21] , \R_DATA_TEMPR9[21] , 
        \R_DATA_TEMPR10[21] , \R_DATA_TEMPR11[21] , 
        \R_DATA_TEMPR12[21] , \R_DATA_TEMPR13[21] , 
        \R_DATA_TEMPR14[21] , \R_DATA_TEMPR15[21] , 
        \R_DATA_TEMPR16[21] , \R_DATA_TEMPR17[21] , 
        \R_DATA_TEMPR18[21] , \R_DATA_TEMPR19[21] , 
        \R_DATA_TEMPR20[21] , \R_DATA_TEMPR21[21] , 
        \R_DATA_TEMPR22[21] , \R_DATA_TEMPR23[21] , 
        \R_DATA_TEMPR24[21] , \R_DATA_TEMPR25[21] , 
        \R_DATA_TEMPR26[21] , \R_DATA_TEMPR27[21] , 
        \R_DATA_TEMPR28[21] , \R_DATA_TEMPR29[21] , 
        \R_DATA_TEMPR30[21] , \R_DATA_TEMPR31[21] , 
        \R_DATA_TEMPR32[21] , \R_DATA_TEMPR33[21] , 
        \R_DATA_TEMPR34[21] , \R_DATA_TEMPR35[21] , 
        \R_DATA_TEMPR36[21] , \R_DATA_TEMPR37[21] , 
        \R_DATA_TEMPR38[21] , \R_DATA_TEMPR39[21] , 
        \R_DATA_TEMPR40[21] , \R_DATA_TEMPR41[21] , 
        \R_DATA_TEMPR42[21] , \R_DATA_TEMPR43[21] , 
        \R_DATA_TEMPR44[21] , \R_DATA_TEMPR45[21] , 
        \R_DATA_TEMPR46[21] , \R_DATA_TEMPR47[21] , 
        \R_DATA_TEMPR48[21] , \R_DATA_TEMPR49[21] , 
        \R_DATA_TEMPR50[21] , \R_DATA_TEMPR51[21] , 
        \R_DATA_TEMPR52[21] , \R_DATA_TEMPR53[21] , 
        \R_DATA_TEMPR54[21] , \R_DATA_TEMPR55[21] , 
        \R_DATA_TEMPR56[21] , \R_DATA_TEMPR57[21] , 
        \R_DATA_TEMPR58[21] , \R_DATA_TEMPR59[21] , 
        \R_DATA_TEMPR60[21] , \R_DATA_TEMPR61[21] , 
        \R_DATA_TEMPR62[21] , \R_DATA_TEMPR63[21] , 
        \R_DATA_TEMPR64[21] , \R_DATA_TEMPR65[21] , 
        \R_DATA_TEMPR66[21] , \R_DATA_TEMPR67[21] , 
        \R_DATA_TEMPR68[21] , \R_DATA_TEMPR69[21] , 
        \R_DATA_TEMPR70[21] , \R_DATA_TEMPR71[21] , 
        \R_DATA_TEMPR72[21] , \R_DATA_TEMPR73[21] , 
        \R_DATA_TEMPR74[21] , \R_DATA_TEMPR75[21] , 
        \R_DATA_TEMPR76[21] , \R_DATA_TEMPR77[21] , 
        \R_DATA_TEMPR78[21] , \R_DATA_TEMPR79[21] , 
        \R_DATA_TEMPR80[21] , \R_DATA_TEMPR81[21] , 
        \R_DATA_TEMPR82[21] , \R_DATA_TEMPR83[21] , 
        \R_DATA_TEMPR84[21] , \R_DATA_TEMPR85[21] , 
        \R_DATA_TEMPR86[21] , \R_DATA_TEMPR87[21] , 
        \R_DATA_TEMPR88[21] , \R_DATA_TEMPR89[21] , 
        \R_DATA_TEMPR90[21] , \R_DATA_TEMPR91[21] , 
        \R_DATA_TEMPR92[21] , \R_DATA_TEMPR93[21] , 
        \R_DATA_TEMPR94[21] , \R_DATA_TEMPR95[21] , 
        \R_DATA_TEMPR96[21] , \R_DATA_TEMPR97[21] , 
        \R_DATA_TEMPR98[21] , \R_DATA_TEMPR99[21] , 
        \R_DATA_TEMPR100[21] , \R_DATA_TEMPR101[21] , 
        \R_DATA_TEMPR102[21] , \R_DATA_TEMPR103[21] , 
        \R_DATA_TEMPR104[21] , \R_DATA_TEMPR105[21] , 
        \R_DATA_TEMPR106[21] , \R_DATA_TEMPR107[21] , 
        \R_DATA_TEMPR108[21] , \R_DATA_TEMPR109[21] , 
        \R_DATA_TEMPR110[21] , \R_DATA_TEMPR111[21] , 
        \R_DATA_TEMPR112[21] , \R_DATA_TEMPR113[21] , 
        \R_DATA_TEMPR114[21] , \R_DATA_TEMPR115[21] , 
        \R_DATA_TEMPR116[21] , \R_DATA_TEMPR117[21] , 
        \R_DATA_TEMPR118[21] , \R_DATA_TEMPR119[21] , 
        \R_DATA_TEMPR120[21] , \R_DATA_TEMPR121[21] , 
        \R_DATA_TEMPR122[21] , \R_DATA_TEMPR123[21] , 
        \R_DATA_TEMPR124[21] , \R_DATA_TEMPR125[21] , 
        \R_DATA_TEMPR126[21] , \R_DATA_TEMPR127[21] , 
        \R_DATA_TEMPR0[22] , \R_DATA_TEMPR1[22] , \R_DATA_TEMPR2[22] , 
        \R_DATA_TEMPR3[22] , \R_DATA_TEMPR4[22] , \R_DATA_TEMPR5[22] , 
        \R_DATA_TEMPR6[22] , \R_DATA_TEMPR7[22] , \R_DATA_TEMPR8[22] , 
        \R_DATA_TEMPR9[22] , \R_DATA_TEMPR10[22] , 
        \R_DATA_TEMPR11[22] , \R_DATA_TEMPR12[22] , 
        \R_DATA_TEMPR13[22] , \R_DATA_TEMPR14[22] , 
        \R_DATA_TEMPR15[22] , \R_DATA_TEMPR16[22] , 
        \R_DATA_TEMPR17[22] , \R_DATA_TEMPR18[22] , 
        \R_DATA_TEMPR19[22] , \R_DATA_TEMPR20[22] , 
        \R_DATA_TEMPR21[22] , \R_DATA_TEMPR22[22] , 
        \R_DATA_TEMPR23[22] , \R_DATA_TEMPR24[22] , 
        \R_DATA_TEMPR25[22] , \R_DATA_TEMPR26[22] , 
        \R_DATA_TEMPR27[22] , \R_DATA_TEMPR28[22] , 
        \R_DATA_TEMPR29[22] , \R_DATA_TEMPR30[22] , 
        \R_DATA_TEMPR31[22] , \R_DATA_TEMPR32[22] , 
        \R_DATA_TEMPR33[22] , \R_DATA_TEMPR34[22] , 
        \R_DATA_TEMPR35[22] , \R_DATA_TEMPR36[22] , 
        \R_DATA_TEMPR37[22] , \R_DATA_TEMPR38[22] , 
        \R_DATA_TEMPR39[22] , \R_DATA_TEMPR40[22] , 
        \R_DATA_TEMPR41[22] , \R_DATA_TEMPR42[22] , 
        \R_DATA_TEMPR43[22] , \R_DATA_TEMPR44[22] , 
        \R_DATA_TEMPR45[22] , \R_DATA_TEMPR46[22] , 
        \R_DATA_TEMPR47[22] , \R_DATA_TEMPR48[22] , 
        \R_DATA_TEMPR49[22] , \R_DATA_TEMPR50[22] , 
        \R_DATA_TEMPR51[22] , \R_DATA_TEMPR52[22] , 
        \R_DATA_TEMPR53[22] , \R_DATA_TEMPR54[22] , 
        \R_DATA_TEMPR55[22] , \R_DATA_TEMPR56[22] , 
        \R_DATA_TEMPR57[22] , \R_DATA_TEMPR58[22] , 
        \R_DATA_TEMPR59[22] , \R_DATA_TEMPR60[22] , 
        \R_DATA_TEMPR61[22] , \R_DATA_TEMPR62[22] , 
        \R_DATA_TEMPR63[22] , \R_DATA_TEMPR64[22] , 
        \R_DATA_TEMPR65[22] , \R_DATA_TEMPR66[22] , 
        \R_DATA_TEMPR67[22] , \R_DATA_TEMPR68[22] , 
        \R_DATA_TEMPR69[22] , \R_DATA_TEMPR70[22] , 
        \R_DATA_TEMPR71[22] , \R_DATA_TEMPR72[22] , 
        \R_DATA_TEMPR73[22] , \R_DATA_TEMPR74[22] , 
        \R_DATA_TEMPR75[22] , \R_DATA_TEMPR76[22] , 
        \R_DATA_TEMPR77[22] , \R_DATA_TEMPR78[22] , 
        \R_DATA_TEMPR79[22] , \R_DATA_TEMPR80[22] , 
        \R_DATA_TEMPR81[22] , \R_DATA_TEMPR82[22] , 
        \R_DATA_TEMPR83[22] , \R_DATA_TEMPR84[22] , 
        \R_DATA_TEMPR85[22] , \R_DATA_TEMPR86[22] , 
        \R_DATA_TEMPR87[22] , \R_DATA_TEMPR88[22] , 
        \R_DATA_TEMPR89[22] , \R_DATA_TEMPR90[22] , 
        \R_DATA_TEMPR91[22] , \R_DATA_TEMPR92[22] , 
        \R_DATA_TEMPR93[22] , \R_DATA_TEMPR94[22] , 
        \R_DATA_TEMPR95[22] , \R_DATA_TEMPR96[22] , 
        \R_DATA_TEMPR97[22] , \R_DATA_TEMPR98[22] , 
        \R_DATA_TEMPR99[22] , \R_DATA_TEMPR100[22] , 
        \R_DATA_TEMPR101[22] , \R_DATA_TEMPR102[22] , 
        \R_DATA_TEMPR103[22] , \R_DATA_TEMPR104[22] , 
        \R_DATA_TEMPR105[22] , \R_DATA_TEMPR106[22] , 
        \R_DATA_TEMPR107[22] , \R_DATA_TEMPR108[22] , 
        \R_DATA_TEMPR109[22] , \R_DATA_TEMPR110[22] , 
        \R_DATA_TEMPR111[22] , \R_DATA_TEMPR112[22] , 
        \R_DATA_TEMPR113[22] , \R_DATA_TEMPR114[22] , 
        \R_DATA_TEMPR115[22] , \R_DATA_TEMPR116[22] , 
        \R_DATA_TEMPR117[22] , \R_DATA_TEMPR118[22] , 
        \R_DATA_TEMPR119[22] , \R_DATA_TEMPR120[22] , 
        \R_DATA_TEMPR121[22] , \R_DATA_TEMPR122[22] , 
        \R_DATA_TEMPR123[22] , \R_DATA_TEMPR124[22] , 
        \R_DATA_TEMPR125[22] , \R_DATA_TEMPR126[22] , 
        \R_DATA_TEMPR127[22] , \R_DATA_TEMPR0[23] , 
        \R_DATA_TEMPR1[23] , \R_DATA_TEMPR2[23] , \R_DATA_TEMPR3[23] , 
        \R_DATA_TEMPR4[23] , \R_DATA_TEMPR5[23] , \R_DATA_TEMPR6[23] , 
        \R_DATA_TEMPR7[23] , \R_DATA_TEMPR8[23] , \R_DATA_TEMPR9[23] , 
        \R_DATA_TEMPR10[23] , \R_DATA_TEMPR11[23] , 
        \R_DATA_TEMPR12[23] , \R_DATA_TEMPR13[23] , 
        \R_DATA_TEMPR14[23] , \R_DATA_TEMPR15[23] , 
        \R_DATA_TEMPR16[23] , \R_DATA_TEMPR17[23] , 
        \R_DATA_TEMPR18[23] , \R_DATA_TEMPR19[23] , 
        \R_DATA_TEMPR20[23] , \R_DATA_TEMPR21[23] , 
        \R_DATA_TEMPR22[23] , \R_DATA_TEMPR23[23] , 
        \R_DATA_TEMPR24[23] , \R_DATA_TEMPR25[23] , 
        \R_DATA_TEMPR26[23] , \R_DATA_TEMPR27[23] , 
        \R_DATA_TEMPR28[23] , \R_DATA_TEMPR29[23] , 
        \R_DATA_TEMPR30[23] , \R_DATA_TEMPR31[23] , 
        \R_DATA_TEMPR32[23] , \R_DATA_TEMPR33[23] , 
        \R_DATA_TEMPR34[23] , \R_DATA_TEMPR35[23] , 
        \R_DATA_TEMPR36[23] , \R_DATA_TEMPR37[23] , 
        \R_DATA_TEMPR38[23] , \R_DATA_TEMPR39[23] , 
        \R_DATA_TEMPR40[23] , \R_DATA_TEMPR41[23] , 
        \R_DATA_TEMPR42[23] , \R_DATA_TEMPR43[23] , 
        \R_DATA_TEMPR44[23] , \R_DATA_TEMPR45[23] , 
        \R_DATA_TEMPR46[23] , \R_DATA_TEMPR47[23] , 
        \R_DATA_TEMPR48[23] , \R_DATA_TEMPR49[23] , 
        \R_DATA_TEMPR50[23] , \R_DATA_TEMPR51[23] , 
        \R_DATA_TEMPR52[23] , \R_DATA_TEMPR53[23] , 
        \R_DATA_TEMPR54[23] , \R_DATA_TEMPR55[23] , 
        \R_DATA_TEMPR56[23] , \R_DATA_TEMPR57[23] , 
        \R_DATA_TEMPR58[23] , \R_DATA_TEMPR59[23] , 
        \R_DATA_TEMPR60[23] , \R_DATA_TEMPR61[23] , 
        \R_DATA_TEMPR62[23] , \R_DATA_TEMPR63[23] , 
        \R_DATA_TEMPR64[23] , \R_DATA_TEMPR65[23] , 
        \R_DATA_TEMPR66[23] , \R_DATA_TEMPR67[23] , 
        \R_DATA_TEMPR68[23] , \R_DATA_TEMPR69[23] , 
        \R_DATA_TEMPR70[23] , \R_DATA_TEMPR71[23] , 
        \R_DATA_TEMPR72[23] , \R_DATA_TEMPR73[23] , 
        \R_DATA_TEMPR74[23] , \R_DATA_TEMPR75[23] , 
        \R_DATA_TEMPR76[23] , \R_DATA_TEMPR77[23] , 
        \R_DATA_TEMPR78[23] , \R_DATA_TEMPR79[23] , 
        \R_DATA_TEMPR80[23] , \R_DATA_TEMPR81[23] , 
        \R_DATA_TEMPR82[23] , \R_DATA_TEMPR83[23] , 
        \R_DATA_TEMPR84[23] , \R_DATA_TEMPR85[23] , 
        \R_DATA_TEMPR86[23] , \R_DATA_TEMPR87[23] , 
        \R_DATA_TEMPR88[23] , \R_DATA_TEMPR89[23] , 
        \R_DATA_TEMPR90[23] , \R_DATA_TEMPR91[23] , 
        \R_DATA_TEMPR92[23] , \R_DATA_TEMPR93[23] , 
        \R_DATA_TEMPR94[23] , \R_DATA_TEMPR95[23] , 
        \R_DATA_TEMPR96[23] , \R_DATA_TEMPR97[23] , 
        \R_DATA_TEMPR98[23] , \R_DATA_TEMPR99[23] , 
        \R_DATA_TEMPR100[23] , \R_DATA_TEMPR101[23] , 
        \R_DATA_TEMPR102[23] , \R_DATA_TEMPR103[23] , 
        \R_DATA_TEMPR104[23] , \R_DATA_TEMPR105[23] , 
        \R_DATA_TEMPR106[23] , \R_DATA_TEMPR107[23] , 
        \R_DATA_TEMPR108[23] , \R_DATA_TEMPR109[23] , 
        \R_DATA_TEMPR110[23] , \R_DATA_TEMPR111[23] , 
        \R_DATA_TEMPR112[23] , \R_DATA_TEMPR113[23] , 
        \R_DATA_TEMPR114[23] , \R_DATA_TEMPR115[23] , 
        \R_DATA_TEMPR116[23] , \R_DATA_TEMPR117[23] , 
        \R_DATA_TEMPR118[23] , \R_DATA_TEMPR119[23] , 
        \R_DATA_TEMPR120[23] , \R_DATA_TEMPR121[23] , 
        \R_DATA_TEMPR122[23] , \R_DATA_TEMPR123[23] , 
        \R_DATA_TEMPR124[23] , \R_DATA_TEMPR125[23] , 
        \R_DATA_TEMPR126[23] , \R_DATA_TEMPR127[23] , 
        \R_DATA_TEMPR0[24] , \R_DATA_TEMPR1[24] , \R_DATA_TEMPR2[24] , 
        \R_DATA_TEMPR3[24] , \R_DATA_TEMPR4[24] , \R_DATA_TEMPR5[24] , 
        \R_DATA_TEMPR6[24] , \R_DATA_TEMPR7[24] , \R_DATA_TEMPR8[24] , 
        \R_DATA_TEMPR9[24] , \R_DATA_TEMPR10[24] , 
        \R_DATA_TEMPR11[24] , \R_DATA_TEMPR12[24] , 
        \R_DATA_TEMPR13[24] , \R_DATA_TEMPR14[24] , 
        \R_DATA_TEMPR15[24] , \R_DATA_TEMPR16[24] , 
        \R_DATA_TEMPR17[24] , \R_DATA_TEMPR18[24] , 
        \R_DATA_TEMPR19[24] , \R_DATA_TEMPR20[24] , 
        \R_DATA_TEMPR21[24] , \R_DATA_TEMPR22[24] , 
        \R_DATA_TEMPR23[24] , \R_DATA_TEMPR24[24] , 
        \R_DATA_TEMPR25[24] , \R_DATA_TEMPR26[24] , 
        \R_DATA_TEMPR27[24] , \R_DATA_TEMPR28[24] , 
        \R_DATA_TEMPR29[24] , \R_DATA_TEMPR30[24] , 
        \R_DATA_TEMPR31[24] , \R_DATA_TEMPR32[24] , 
        \R_DATA_TEMPR33[24] , \R_DATA_TEMPR34[24] , 
        \R_DATA_TEMPR35[24] , \R_DATA_TEMPR36[24] , 
        \R_DATA_TEMPR37[24] , \R_DATA_TEMPR38[24] , 
        \R_DATA_TEMPR39[24] , \R_DATA_TEMPR40[24] , 
        \R_DATA_TEMPR41[24] , \R_DATA_TEMPR42[24] , 
        \R_DATA_TEMPR43[24] , \R_DATA_TEMPR44[24] , 
        \R_DATA_TEMPR45[24] , \R_DATA_TEMPR46[24] , 
        \R_DATA_TEMPR47[24] , \R_DATA_TEMPR48[24] , 
        \R_DATA_TEMPR49[24] , \R_DATA_TEMPR50[24] , 
        \R_DATA_TEMPR51[24] , \R_DATA_TEMPR52[24] , 
        \R_DATA_TEMPR53[24] , \R_DATA_TEMPR54[24] , 
        \R_DATA_TEMPR55[24] , \R_DATA_TEMPR56[24] , 
        \R_DATA_TEMPR57[24] , \R_DATA_TEMPR58[24] , 
        \R_DATA_TEMPR59[24] , \R_DATA_TEMPR60[24] , 
        \R_DATA_TEMPR61[24] , \R_DATA_TEMPR62[24] , 
        \R_DATA_TEMPR63[24] , \R_DATA_TEMPR64[24] , 
        \R_DATA_TEMPR65[24] , \R_DATA_TEMPR66[24] , 
        \R_DATA_TEMPR67[24] , \R_DATA_TEMPR68[24] , 
        \R_DATA_TEMPR69[24] , \R_DATA_TEMPR70[24] , 
        \R_DATA_TEMPR71[24] , \R_DATA_TEMPR72[24] , 
        \R_DATA_TEMPR73[24] , \R_DATA_TEMPR74[24] , 
        \R_DATA_TEMPR75[24] , \R_DATA_TEMPR76[24] , 
        \R_DATA_TEMPR77[24] , \R_DATA_TEMPR78[24] , 
        \R_DATA_TEMPR79[24] , \R_DATA_TEMPR80[24] , 
        \R_DATA_TEMPR81[24] , \R_DATA_TEMPR82[24] , 
        \R_DATA_TEMPR83[24] , \R_DATA_TEMPR84[24] , 
        \R_DATA_TEMPR85[24] , \R_DATA_TEMPR86[24] , 
        \R_DATA_TEMPR87[24] , \R_DATA_TEMPR88[24] , 
        \R_DATA_TEMPR89[24] , \R_DATA_TEMPR90[24] , 
        \R_DATA_TEMPR91[24] , \R_DATA_TEMPR92[24] , 
        \R_DATA_TEMPR93[24] , \R_DATA_TEMPR94[24] , 
        \R_DATA_TEMPR95[24] , \R_DATA_TEMPR96[24] , 
        \R_DATA_TEMPR97[24] , \R_DATA_TEMPR98[24] , 
        \R_DATA_TEMPR99[24] , \R_DATA_TEMPR100[24] , 
        \R_DATA_TEMPR101[24] , \R_DATA_TEMPR102[24] , 
        \R_DATA_TEMPR103[24] , \R_DATA_TEMPR104[24] , 
        \R_DATA_TEMPR105[24] , \R_DATA_TEMPR106[24] , 
        \R_DATA_TEMPR107[24] , \R_DATA_TEMPR108[24] , 
        \R_DATA_TEMPR109[24] , \R_DATA_TEMPR110[24] , 
        \R_DATA_TEMPR111[24] , \R_DATA_TEMPR112[24] , 
        \R_DATA_TEMPR113[24] , \R_DATA_TEMPR114[24] , 
        \R_DATA_TEMPR115[24] , \R_DATA_TEMPR116[24] , 
        \R_DATA_TEMPR117[24] , \R_DATA_TEMPR118[24] , 
        \R_DATA_TEMPR119[24] , \R_DATA_TEMPR120[24] , 
        \R_DATA_TEMPR121[24] , \R_DATA_TEMPR122[24] , 
        \R_DATA_TEMPR123[24] , \R_DATA_TEMPR124[24] , 
        \R_DATA_TEMPR125[24] , \R_DATA_TEMPR126[24] , 
        \R_DATA_TEMPR127[24] , \R_DATA_TEMPR0[25] , 
        \R_DATA_TEMPR1[25] , \R_DATA_TEMPR2[25] , \R_DATA_TEMPR3[25] , 
        \R_DATA_TEMPR4[25] , \R_DATA_TEMPR5[25] , \R_DATA_TEMPR6[25] , 
        \R_DATA_TEMPR7[25] , \R_DATA_TEMPR8[25] , \R_DATA_TEMPR9[25] , 
        \R_DATA_TEMPR10[25] , \R_DATA_TEMPR11[25] , 
        \R_DATA_TEMPR12[25] , \R_DATA_TEMPR13[25] , 
        \R_DATA_TEMPR14[25] , \R_DATA_TEMPR15[25] , 
        \R_DATA_TEMPR16[25] , \R_DATA_TEMPR17[25] , 
        \R_DATA_TEMPR18[25] , \R_DATA_TEMPR19[25] , 
        \R_DATA_TEMPR20[25] , \R_DATA_TEMPR21[25] , 
        \R_DATA_TEMPR22[25] , \R_DATA_TEMPR23[25] , 
        \R_DATA_TEMPR24[25] , \R_DATA_TEMPR25[25] , 
        \R_DATA_TEMPR26[25] , \R_DATA_TEMPR27[25] , 
        \R_DATA_TEMPR28[25] , \R_DATA_TEMPR29[25] , 
        \R_DATA_TEMPR30[25] , \R_DATA_TEMPR31[25] , 
        \R_DATA_TEMPR32[25] , \R_DATA_TEMPR33[25] , 
        \R_DATA_TEMPR34[25] , \R_DATA_TEMPR35[25] , 
        \R_DATA_TEMPR36[25] , \R_DATA_TEMPR37[25] , 
        \R_DATA_TEMPR38[25] , \R_DATA_TEMPR39[25] , 
        \R_DATA_TEMPR40[25] , \R_DATA_TEMPR41[25] , 
        \R_DATA_TEMPR42[25] , \R_DATA_TEMPR43[25] , 
        \R_DATA_TEMPR44[25] , \R_DATA_TEMPR45[25] , 
        \R_DATA_TEMPR46[25] , \R_DATA_TEMPR47[25] , 
        \R_DATA_TEMPR48[25] , \R_DATA_TEMPR49[25] , 
        \R_DATA_TEMPR50[25] , \R_DATA_TEMPR51[25] , 
        \R_DATA_TEMPR52[25] , \R_DATA_TEMPR53[25] , 
        \R_DATA_TEMPR54[25] , \R_DATA_TEMPR55[25] , 
        \R_DATA_TEMPR56[25] , \R_DATA_TEMPR57[25] , 
        \R_DATA_TEMPR58[25] , \R_DATA_TEMPR59[25] , 
        \R_DATA_TEMPR60[25] , \R_DATA_TEMPR61[25] , 
        \R_DATA_TEMPR62[25] , \R_DATA_TEMPR63[25] , 
        \R_DATA_TEMPR64[25] , \R_DATA_TEMPR65[25] , 
        \R_DATA_TEMPR66[25] , \R_DATA_TEMPR67[25] , 
        \R_DATA_TEMPR68[25] , \R_DATA_TEMPR69[25] , 
        \R_DATA_TEMPR70[25] , \R_DATA_TEMPR71[25] , 
        \R_DATA_TEMPR72[25] , \R_DATA_TEMPR73[25] , 
        \R_DATA_TEMPR74[25] , \R_DATA_TEMPR75[25] , 
        \R_DATA_TEMPR76[25] , \R_DATA_TEMPR77[25] , 
        \R_DATA_TEMPR78[25] , \R_DATA_TEMPR79[25] , 
        \R_DATA_TEMPR80[25] , \R_DATA_TEMPR81[25] , 
        \R_DATA_TEMPR82[25] , \R_DATA_TEMPR83[25] , 
        \R_DATA_TEMPR84[25] , \R_DATA_TEMPR85[25] , 
        \R_DATA_TEMPR86[25] , \R_DATA_TEMPR87[25] , 
        \R_DATA_TEMPR88[25] , \R_DATA_TEMPR89[25] , 
        \R_DATA_TEMPR90[25] , \R_DATA_TEMPR91[25] , 
        \R_DATA_TEMPR92[25] , \R_DATA_TEMPR93[25] , 
        \R_DATA_TEMPR94[25] , \R_DATA_TEMPR95[25] , 
        \R_DATA_TEMPR96[25] , \R_DATA_TEMPR97[25] , 
        \R_DATA_TEMPR98[25] , \R_DATA_TEMPR99[25] , 
        \R_DATA_TEMPR100[25] , \R_DATA_TEMPR101[25] , 
        \R_DATA_TEMPR102[25] , \R_DATA_TEMPR103[25] , 
        \R_DATA_TEMPR104[25] , \R_DATA_TEMPR105[25] , 
        \R_DATA_TEMPR106[25] , \R_DATA_TEMPR107[25] , 
        \R_DATA_TEMPR108[25] , \R_DATA_TEMPR109[25] , 
        \R_DATA_TEMPR110[25] , \R_DATA_TEMPR111[25] , 
        \R_DATA_TEMPR112[25] , \R_DATA_TEMPR113[25] , 
        \R_DATA_TEMPR114[25] , \R_DATA_TEMPR115[25] , 
        \R_DATA_TEMPR116[25] , \R_DATA_TEMPR117[25] , 
        \R_DATA_TEMPR118[25] , \R_DATA_TEMPR119[25] , 
        \R_DATA_TEMPR120[25] , \R_DATA_TEMPR121[25] , 
        \R_DATA_TEMPR122[25] , \R_DATA_TEMPR123[25] , 
        \R_DATA_TEMPR124[25] , \R_DATA_TEMPR125[25] , 
        \R_DATA_TEMPR126[25] , \R_DATA_TEMPR127[25] , 
        \R_DATA_TEMPR0[26] , \R_DATA_TEMPR1[26] , \R_DATA_TEMPR2[26] , 
        \R_DATA_TEMPR3[26] , \R_DATA_TEMPR4[26] , \R_DATA_TEMPR5[26] , 
        \R_DATA_TEMPR6[26] , \R_DATA_TEMPR7[26] , \R_DATA_TEMPR8[26] , 
        \R_DATA_TEMPR9[26] , \R_DATA_TEMPR10[26] , 
        \R_DATA_TEMPR11[26] , \R_DATA_TEMPR12[26] , 
        \R_DATA_TEMPR13[26] , \R_DATA_TEMPR14[26] , 
        \R_DATA_TEMPR15[26] , \R_DATA_TEMPR16[26] , 
        \R_DATA_TEMPR17[26] , \R_DATA_TEMPR18[26] , 
        \R_DATA_TEMPR19[26] , \R_DATA_TEMPR20[26] , 
        \R_DATA_TEMPR21[26] , \R_DATA_TEMPR22[26] , 
        \R_DATA_TEMPR23[26] , \R_DATA_TEMPR24[26] , 
        \R_DATA_TEMPR25[26] , \R_DATA_TEMPR26[26] , 
        \R_DATA_TEMPR27[26] , \R_DATA_TEMPR28[26] , 
        \R_DATA_TEMPR29[26] , \R_DATA_TEMPR30[26] , 
        \R_DATA_TEMPR31[26] , \R_DATA_TEMPR32[26] , 
        \R_DATA_TEMPR33[26] , \R_DATA_TEMPR34[26] , 
        \R_DATA_TEMPR35[26] , \R_DATA_TEMPR36[26] , 
        \R_DATA_TEMPR37[26] , \R_DATA_TEMPR38[26] , 
        \R_DATA_TEMPR39[26] , \R_DATA_TEMPR40[26] , 
        \R_DATA_TEMPR41[26] , \R_DATA_TEMPR42[26] , 
        \R_DATA_TEMPR43[26] , \R_DATA_TEMPR44[26] , 
        \R_DATA_TEMPR45[26] , \R_DATA_TEMPR46[26] , 
        \R_DATA_TEMPR47[26] , \R_DATA_TEMPR48[26] , 
        \R_DATA_TEMPR49[26] , \R_DATA_TEMPR50[26] , 
        \R_DATA_TEMPR51[26] , \R_DATA_TEMPR52[26] , 
        \R_DATA_TEMPR53[26] , \R_DATA_TEMPR54[26] , 
        \R_DATA_TEMPR55[26] , \R_DATA_TEMPR56[26] , 
        \R_DATA_TEMPR57[26] , \R_DATA_TEMPR58[26] , 
        \R_DATA_TEMPR59[26] , \R_DATA_TEMPR60[26] , 
        \R_DATA_TEMPR61[26] , \R_DATA_TEMPR62[26] , 
        \R_DATA_TEMPR63[26] , \R_DATA_TEMPR64[26] , 
        \R_DATA_TEMPR65[26] , \R_DATA_TEMPR66[26] , 
        \R_DATA_TEMPR67[26] , \R_DATA_TEMPR68[26] , 
        \R_DATA_TEMPR69[26] , \R_DATA_TEMPR70[26] , 
        \R_DATA_TEMPR71[26] , \R_DATA_TEMPR72[26] , 
        \R_DATA_TEMPR73[26] , \R_DATA_TEMPR74[26] , 
        \R_DATA_TEMPR75[26] , \R_DATA_TEMPR76[26] , 
        \R_DATA_TEMPR77[26] , \R_DATA_TEMPR78[26] , 
        \R_DATA_TEMPR79[26] , \R_DATA_TEMPR80[26] , 
        \R_DATA_TEMPR81[26] , \R_DATA_TEMPR82[26] , 
        \R_DATA_TEMPR83[26] , \R_DATA_TEMPR84[26] , 
        \R_DATA_TEMPR85[26] , \R_DATA_TEMPR86[26] , 
        \R_DATA_TEMPR87[26] , \R_DATA_TEMPR88[26] , 
        \R_DATA_TEMPR89[26] , \R_DATA_TEMPR90[26] , 
        \R_DATA_TEMPR91[26] , \R_DATA_TEMPR92[26] , 
        \R_DATA_TEMPR93[26] , \R_DATA_TEMPR94[26] , 
        \R_DATA_TEMPR95[26] , \R_DATA_TEMPR96[26] , 
        \R_DATA_TEMPR97[26] , \R_DATA_TEMPR98[26] , 
        \R_DATA_TEMPR99[26] , \R_DATA_TEMPR100[26] , 
        \R_DATA_TEMPR101[26] , \R_DATA_TEMPR102[26] , 
        \R_DATA_TEMPR103[26] , \R_DATA_TEMPR104[26] , 
        \R_DATA_TEMPR105[26] , \R_DATA_TEMPR106[26] , 
        \R_DATA_TEMPR107[26] , \R_DATA_TEMPR108[26] , 
        \R_DATA_TEMPR109[26] , \R_DATA_TEMPR110[26] , 
        \R_DATA_TEMPR111[26] , \R_DATA_TEMPR112[26] , 
        \R_DATA_TEMPR113[26] , \R_DATA_TEMPR114[26] , 
        \R_DATA_TEMPR115[26] , \R_DATA_TEMPR116[26] , 
        \R_DATA_TEMPR117[26] , \R_DATA_TEMPR118[26] , 
        \R_DATA_TEMPR119[26] , \R_DATA_TEMPR120[26] , 
        \R_DATA_TEMPR121[26] , \R_DATA_TEMPR122[26] , 
        \R_DATA_TEMPR123[26] , \R_DATA_TEMPR124[26] , 
        \R_DATA_TEMPR125[26] , \R_DATA_TEMPR126[26] , 
        \R_DATA_TEMPR127[26] , \R_DATA_TEMPR0[27] , 
        \R_DATA_TEMPR1[27] , \R_DATA_TEMPR2[27] , \R_DATA_TEMPR3[27] , 
        \R_DATA_TEMPR4[27] , \R_DATA_TEMPR5[27] , \R_DATA_TEMPR6[27] , 
        \R_DATA_TEMPR7[27] , \R_DATA_TEMPR8[27] , \R_DATA_TEMPR9[27] , 
        \R_DATA_TEMPR10[27] , \R_DATA_TEMPR11[27] , 
        \R_DATA_TEMPR12[27] , \R_DATA_TEMPR13[27] , 
        \R_DATA_TEMPR14[27] , \R_DATA_TEMPR15[27] , 
        \R_DATA_TEMPR16[27] , \R_DATA_TEMPR17[27] , 
        \R_DATA_TEMPR18[27] , \R_DATA_TEMPR19[27] , 
        \R_DATA_TEMPR20[27] , \R_DATA_TEMPR21[27] , 
        \R_DATA_TEMPR22[27] , \R_DATA_TEMPR23[27] , 
        \R_DATA_TEMPR24[27] , \R_DATA_TEMPR25[27] , 
        \R_DATA_TEMPR26[27] , \R_DATA_TEMPR27[27] , 
        \R_DATA_TEMPR28[27] , \R_DATA_TEMPR29[27] , 
        \R_DATA_TEMPR30[27] , \R_DATA_TEMPR31[27] , 
        \R_DATA_TEMPR32[27] , \R_DATA_TEMPR33[27] , 
        \R_DATA_TEMPR34[27] , \R_DATA_TEMPR35[27] , 
        \R_DATA_TEMPR36[27] , \R_DATA_TEMPR37[27] , 
        \R_DATA_TEMPR38[27] , \R_DATA_TEMPR39[27] , 
        \R_DATA_TEMPR40[27] , \R_DATA_TEMPR41[27] , 
        \R_DATA_TEMPR42[27] , \R_DATA_TEMPR43[27] , 
        \R_DATA_TEMPR44[27] , \R_DATA_TEMPR45[27] , 
        \R_DATA_TEMPR46[27] , \R_DATA_TEMPR47[27] , 
        \R_DATA_TEMPR48[27] , \R_DATA_TEMPR49[27] , 
        \R_DATA_TEMPR50[27] , \R_DATA_TEMPR51[27] , 
        \R_DATA_TEMPR52[27] , \R_DATA_TEMPR53[27] , 
        \R_DATA_TEMPR54[27] , \R_DATA_TEMPR55[27] , 
        \R_DATA_TEMPR56[27] , \R_DATA_TEMPR57[27] , 
        \R_DATA_TEMPR58[27] , \R_DATA_TEMPR59[27] , 
        \R_DATA_TEMPR60[27] , \R_DATA_TEMPR61[27] , 
        \R_DATA_TEMPR62[27] , \R_DATA_TEMPR63[27] , 
        \R_DATA_TEMPR64[27] , \R_DATA_TEMPR65[27] , 
        \R_DATA_TEMPR66[27] , \R_DATA_TEMPR67[27] , 
        \R_DATA_TEMPR68[27] , \R_DATA_TEMPR69[27] , 
        \R_DATA_TEMPR70[27] , \R_DATA_TEMPR71[27] , 
        \R_DATA_TEMPR72[27] , \R_DATA_TEMPR73[27] , 
        \R_DATA_TEMPR74[27] , \R_DATA_TEMPR75[27] , 
        \R_DATA_TEMPR76[27] , \R_DATA_TEMPR77[27] , 
        \R_DATA_TEMPR78[27] , \R_DATA_TEMPR79[27] , 
        \R_DATA_TEMPR80[27] , \R_DATA_TEMPR81[27] , 
        \R_DATA_TEMPR82[27] , \R_DATA_TEMPR83[27] , 
        \R_DATA_TEMPR84[27] , \R_DATA_TEMPR85[27] , 
        \R_DATA_TEMPR86[27] , \R_DATA_TEMPR87[27] , 
        \R_DATA_TEMPR88[27] , \R_DATA_TEMPR89[27] , 
        \R_DATA_TEMPR90[27] , \R_DATA_TEMPR91[27] , 
        \R_DATA_TEMPR92[27] , \R_DATA_TEMPR93[27] , 
        \R_DATA_TEMPR94[27] , \R_DATA_TEMPR95[27] , 
        \R_DATA_TEMPR96[27] , \R_DATA_TEMPR97[27] , 
        \R_DATA_TEMPR98[27] , \R_DATA_TEMPR99[27] , 
        \R_DATA_TEMPR100[27] , \R_DATA_TEMPR101[27] , 
        \R_DATA_TEMPR102[27] , \R_DATA_TEMPR103[27] , 
        \R_DATA_TEMPR104[27] , \R_DATA_TEMPR105[27] , 
        \R_DATA_TEMPR106[27] , \R_DATA_TEMPR107[27] , 
        \R_DATA_TEMPR108[27] , \R_DATA_TEMPR109[27] , 
        \R_DATA_TEMPR110[27] , \R_DATA_TEMPR111[27] , 
        \R_DATA_TEMPR112[27] , \R_DATA_TEMPR113[27] , 
        \R_DATA_TEMPR114[27] , \R_DATA_TEMPR115[27] , 
        \R_DATA_TEMPR116[27] , \R_DATA_TEMPR117[27] , 
        \R_DATA_TEMPR118[27] , \R_DATA_TEMPR119[27] , 
        \R_DATA_TEMPR120[27] , \R_DATA_TEMPR121[27] , 
        \R_DATA_TEMPR122[27] , \R_DATA_TEMPR123[27] , 
        \R_DATA_TEMPR124[27] , \R_DATA_TEMPR125[27] , 
        \R_DATA_TEMPR126[27] , \R_DATA_TEMPR127[27] , 
        \R_DATA_TEMPR0[28] , \R_DATA_TEMPR1[28] , \R_DATA_TEMPR2[28] , 
        \R_DATA_TEMPR3[28] , \R_DATA_TEMPR4[28] , \R_DATA_TEMPR5[28] , 
        \R_DATA_TEMPR6[28] , \R_DATA_TEMPR7[28] , \R_DATA_TEMPR8[28] , 
        \R_DATA_TEMPR9[28] , \R_DATA_TEMPR10[28] , 
        \R_DATA_TEMPR11[28] , \R_DATA_TEMPR12[28] , 
        \R_DATA_TEMPR13[28] , \R_DATA_TEMPR14[28] , 
        \R_DATA_TEMPR15[28] , \R_DATA_TEMPR16[28] , 
        \R_DATA_TEMPR17[28] , \R_DATA_TEMPR18[28] , 
        \R_DATA_TEMPR19[28] , \R_DATA_TEMPR20[28] , 
        \R_DATA_TEMPR21[28] , \R_DATA_TEMPR22[28] , 
        \R_DATA_TEMPR23[28] , \R_DATA_TEMPR24[28] , 
        \R_DATA_TEMPR25[28] , \R_DATA_TEMPR26[28] , 
        \R_DATA_TEMPR27[28] , \R_DATA_TEMPR28[28] , 
        \R_DATA_TEMPR29[28] , \R_DATA_TEMPR30[28] , 
        \R_DATA_TEMPR31[28] , \R_DATA_TEMPR32[28] , 
        \R_DATA_TEMPR33[28] , \R_DATA_TEMPR34[28] , 
        \R_DATA_TEMPR35[28] , \R_DATA_TEMPR36[28] , 
        \R_DATA_TEMPR37[28] , \R_DATA_TEMPR38[28] , 
        \R_DATA_TEMPR39[28] , \R_DATA_TEMPR40[28] , 
        \R_DATA_TEMPR41[28] , \R_DATA_TEMPR42[28] , 
        \R_DATA_TEMPR43[28] , \R_DATA_TEMPR44[28] , 
        \R_DATA_TEMPR45[28] , \R_DATA_TEMPR46[28] , 
        \R_DATA_TEMPR47[28] , \R_DATA_TEMPR48[28] , 
        \R_DATA_TEMPR49[28] , \R_DATA_TEMPR50[28] , 
        \R_DATA_TEMPR51[28] , \R_DATA_TEMPR52[28] , 
        \R_DATA_TEMPR53[28] , \R_DATA_TEMPR54[28] , 
        \R_DATA_TEMPR55[28] , \R_DATA_TEMPR56[28] , 
        \R_DATA_TEMPR57[28] , \R_DATA_TEMPR58[28] , 
        \R_DATA_TEMPR59[28] , \R_DATA_TEMPR60[28] , 
        \R_DATA_TEMPR61[28] , \R_DATA_TEMPR62[28] , 
        \R_DATA_TEMPR63[28] , \R_DATA_TEMPR64[28] , 
        \R_DATA_TEMPR65[28] , \R_DATA_TEMPR66[28] , 
        \R_DATA_TEMPR67[28] , \R_DATA_TEMPR68[28] , 
        \R_DATA_TEMPR69[28] , \R_DATA_TEMPR70[28] , 
        \R_DATA_TEMPR71[28] , \R_DATA_TEMPR72[28] , 
        \R_DATA_TEMPR73[28] , \R_DATA_TEMPR74[28] , 
        \R_DATA_TEMPR75[28] , \R_DATA_TEMPR76[28] , 
        \R_DATA_TEMPR77[28] , \R_DATA_TEMPR78[28] , 
        \R_DATA_TEMPR79[28] , \R_DATA_TEMPR80[28] , 
        \R_DATA_TEMPR81[28] , \R_DATA_TEMPR82[28] , 
        \R_DATA_TEMPR83[28] , \R_DATA_TEMPR84[28] , 
        \R_DATA_TEMPR85[28] , \R_DATA_TEMPR86[28] , 
        \R_DATA_TEMPR87[28] , \R_DATA_TEMPR88[28] , 
        \R_DATA_TEMPR89[28] , \R_DATA_TEMPR90[28] , 
        \R_DATA_TEMPR91[28] , \R_DATA_TEMPR92[28] , 
        \R_DATA_TEMPR93[28] , \R_DATA_TEMPR94[28] , 
        \R_DATA_TEMPR95[28] , \R_DATA_TEMPR96[28] , 
        \R_DATA_TEMPR97[28] , \R_DATA_TEMPR98[28] , 
        \R_DATA_TEMPR99[28] , \R_DATA_TEMPR100[28] , 
        \R_DATA_TEMPR101[28] , \R_DATA_TEMPR102[28] , 
        \R_DATA_TEMPR103[28] , \R_DATA_TEMPR104[28] , 
        \R_DATA_TEMPR105[28] , \R_DATA_TEMPR106[28] , 
        \R_DATA_TEMPR107[28] , \R_DATA_TEMPR108[28] , 
        \R_DATA_TEMPR109[28] , \R_DATA_TEMPR110[28] , 
        \R_DATA_TEMPR111[28] , \R_DATA_TEMPR112[28] , 
        \R_DATA_TEMPR113[28] , \R_DATA_TEMPR114[28] , 
        \R_DATA_TEMPR115[28] , \R_DATA_TEMPR116[28] , 
        \R_DATA_TEMPR117[28] , \R_DATA_TEMPR118[28] , 
        \R_DATA_TEMPR119[28] , \R_DATA_TEMPR120[28] , 
        \R_DATA_TEMPR121[28] , \R_DATA_TEMPR122[28] , 
        \R_DATA_TEMPR123[28] , \R_DATA_TEMPR124[28] , 
        \R_DATA_TEMPR125[28] , \R_DATA_TEMPR126[28] , 
        \R_DATA_TEMPR127[28] , \R_DATA_TEMPR0[29] , 
        \R_DATA_TEMPR1[29] , \R_DATA_TEMPR2[29] , \R_DATA_TEMPR3[29] , 
        \R_DATA_TEMPR4[29] , \R_DATA_TEMPR5[29] , \R_DATA_TEMPR6[29] , 
        \R_DATA_TEMPR7[29] , \R_DATA_TEMPR8[29] , \R_DATA_TEMPR9[29] , 
        \R_DATA_TEMPR10[29] , \R_DATA_TEMPR11[29] , 
        \R_DATA_TEMPR12[29] , \R_DATA_TEMPR13[29] , 
        \R_DATA_TEMPR14[29] , \R_DATA_TEMPR15[29] , 
        \R_DATA_TEMPR16[29] , \R_DATA_TEMPR17[29] , 
        \R_DATA_TEMPR18[29] , \R_DATA_TEMPR19[29] , 
        \R_DATA_TEMPR20[29] , \R_DATA_TEMPR21[29] , 
        \R_DATA_TEMPR22[29] , \R_DATA_TEMPR23[29] , 
        \R_DATA_TEMPR24[29] , \R_DATA_TEMPR25[29] , 
        \R_DATA_TEMPR26[29] , \R_DATA_TEMPR27[29] , 
        \R_DATA_TEMPR28[29] , \R_DATA_TEMPR29[29] , 
        \R_DATA_TEMPR30[29] , \R_DATA_TEMPR31[29] , 
        \R_DATA_TEMPR32[29] , \R_DATA_TEMPR33[29] , 
        \R_DATA_TEMPR34[29] , \R_DATA_TEMPR35[29] , 
        \R_DATA_TEMPR36[29] , \R_DATA_TEMPR37[29] , 
        \R_DATA_TEMPR38[29] , \R_DATA_TEMPR39[29] , 
        \R_DATA_TEMPR40[29] , \R_DATA_TEMPR41[29] , 
        \R_DATA_TEMPR42[29] , \R_DATA_TEMPR43[29] , 
        \R_DATA_TEMPR44[29] , \R_DATA_TEMPR45[29] , 
        \R_DATA_TEMPR46[29] , \R_DATA_TEMPR47[29] , 
        \R_DATA_TEMPR48[29] , \R_DATA_TEMPR49[29] , 
        \R_DATA_TEMPR50[29] , \R_DATA_TEMPR51[29] , 
        \R_DATA_TEMPR52[29] , \R_DATA_TEMPR53[29] , 
        \R_DATA_TEMPR54[29] , \R_DATA_TEMPR55[29] , 
        \R_DATA_TEMPR56[29] , \R_DATA_TEMPR57[29] , 
        \R_DATA_TEMPR58[29] , \R_DATA_TEMPR59[29] , 
        \R_DATA_TEMPR60[29] , \R_DATA_TEMPR61[29] , 
        \R_DATA_TEMPR62[29] , \R_DATA_TEMPR63[29] , 
        \R_DATA_TEMPR64[29] , \R_DATA_TEMPR65[29] , 
        \R_DATA_TEMPR66[29] , \R_DATA_TEMPR67[29] , 
        \R_DATA_TEMPR68[29] , \R_DATA_TEMPR69[29] , 
        \R_DATA_TEMPR70[29] , \R_DATA_TEMPR71[29] , 
        \R_DATA_TEMPR72[29] , \R_DATA_TEMPR73[29] , 
        \R_DATA_TEMPR74[29] , \R_DATA_TEMPR75[29] , 
        \R_DATA_TEMPR76[29] , \R_DATA_TEMPR77[29] , 
        \R_DATA_TEMPR78[29] , \R_DATA_TEMPR79[29] , 
        \R_DATA_TEMPR80[29] , \R_DATA_TEMPR81[29] , 
        \R_DATA_TEMPR82[29] , \R_DATA_TEMPR83[29] , 
        \R_DATA_TEMPR84[29] , \R_DATA_TEMPR85[29] , 
        \R_DATA_TEMPR86[29] , \R_DATA_TEMPR87[29] , 
        \R_DATA_TEMPR88[29] , \R_DATA_TEMPR89[29] , 
        \R_DATA_TEMPR90[29] , \R_DATA_TEMPR91[29] , 
        \R_DATA_TEMPR92[29] , \R_DATA_TEMPR93[29] , 
        \R_DATA_TEMPR94[29] , \R_DATA_TEMPR95[29] , 
        \R_DATA_TEMPR96[29] , \R_DATA_TEMPR97[29] , 
        \R_DATA_TEMPR98[29] , \R_DATA_TEMPR99[29] , 
        \R_DATA_TEMPR100[29] , \R_DATA_TEMPR101[29] , 
        \R_DATA_TEMPR102[29] , \R_DATA_TEMPR103[29] , 
        \R_DATA_TEMPR104[29] , \R_DATA_TEMPR105[29] , 
        \R_DATA_TEMPR106[29] , \R_DATA_TEMPR107[29] , 
        \R_DATA_TEMPR108[29] , \R_DATA_TEMPR109[29] , 
        \R_DATA_TEMPR110[29] , \R_DATA_TEMPR111[29] , 
        \R_DATA_TEMPR112[29] , \R_DATA_TEMPR113[29] , 
        \R_DATA_TEMPR114[29] , \R_DATA_TEMPR115[29] , 
        \R_DATA_TEMPR116[29] , \R_DATA_TEMPR117[29] , 
        \R_DATA_TEMPR118[29] , \R_DATA_TEMPR119[29] , 
        \R_DATA_TEMPR120[29] , \R_DATA_TEMPR121[29] , 
        \R_DATA_TEMPR122[29] , \R_DATA_TEMPR123[29] , 
        \R_DATA_TEMPR124[29] , \R_DATA_TEMPR125[29] , 
        \R_DATA_TEMPR126[29] , \R_DATA_TEMPR127[29] , 
        \R_DATA_TEMPR0[30] , \R_DATA_TEMPR1[30] , \R_DATA_TEMPR2[30] , 
        \R_DATA_TEMPR3[30] , \R_DATA_TEMPR4[30] , \R_DATA_TEMPR5[30] , 
        \R_DATA_TEMPR6[30] , \R_DATA_TEMPR7[30] , \R_DATA_TEMPR8[30] , 
        \R_DATA_TEMPR9[30] , \R_DATA_TEMPR10[30] , 
        \R_DATA_TEMPR11[30] , \R_DATA_TEMPR12[30] , 
        \R_DATA_TEMPR13[30] , \R_DATA_TEMPR14[30] , 
        \R_DATA_TEMPR15[30] , \R_DATA_TEMPR16[30] , 
        \R_DATA_TEMPR17[30] , \R_DATA_TEMPR18[30] , 
        \R_DATA_TEMPR19[30] , \R_DATA_TEMPR20[30] , 
        \R_DATA_TEMPR21[30] , \R_DATA_TEMPR22[30] , 
        \R_DATA_TEMPR23[30] , \R_DATA_TEMPR24[30] , 
        \R_DATA_TEMPR25[30] , \R_DATA_TEMPR26[30] , 
        \R_DATA_TEMPR27[30] , \R_DATA_TEMPR28[30] , 
        \R_DATA_TEMPR29[30] , \R_DATA_TEMPR30[30] , 
        \R_DATA_TEMPR31[30] , \R_DATA_TEMPR32[30] , 
        \R_DATA_TEMPR33[30] , \R_DATA_TEMPR34[30] , 
        \R_DATA_TEMPR35[30] , \R_DATA_TEMPR36[30] , 
        \R_DATA_TEMPR37[30] , \R_DATA_TEMPR38[30] , 
        \R_DATA_TEMPR39[30] , \R_DATA_TEMPR40[30] , 
        \R_DATA_TEMPR41[30] , \R_DATA_TEMPR42[30] , 
        \R_DATA_TEMPR43[30] , \R_DATA_TEMPR44[30] , 
        \R_DATA_TEMPR45[30] , \R_DATA_TEMPR46[30] , 
        \R_DATA_TEMPR47[30] , \R_DATA_TEMPR48[30] , 
        \R_DATA_TEMPR49[30] , \R_DATA_TEMPR50[30] , 
        \R_DATA_TEMPR51[30] , \R_DATA_TEMPR52[30] , 
        \R_DATA_TEMPR53[30] , \R_DATA_TEMPR54[30] , 
        \R_DATA_TEMPR55[30] , \R_DATA_TEMPR56[30] , 
        \R_DATA_TEMPR57[30] , \R_DATA_TEMPR58[30] , 
        \R_DATA_TEMPR59[30] , \R_DATA_TEMPR60[30] , 
        \R_DATA_TEMPR61[30] , \R_DATA_TEMPR62[30] , 
        \R_DATA_TEMPR63[30] , \R_DATA_TEMPR64[30] , 
        \R_DATA_TEMPR65[30] , \R_DATA_TEMPR66[30] , 
        \R_DATA_TEMPR67[30] , \R_DATA_TEMPR68[30] , 
        \R_DATA_TEMPR69[30] , \R_DATA_TEMPR70[30] , 
        \R_DATA_TEMPR71[30] , \R_DATA_TEMPR72[30] , 
        \R_DATA_TEMPR73[30] , \R_DATA_TEMPR74[30] , 
        \R_DATA_TEMPR75[30] , \R_DATA_TEMPR76[30] , 
        \R_DATA_TEMPR77[30] , \R_DATA_TEMPR78[30] , 
        \R_DATA_TEMPR79[30] , \R_DATA_TEMPR80[30] , 
        \R_DATA_TEMPR81[30] , \R_DATA_TEMPR82[30] , 
        \R_DATA_TEMPR83[30] , \R_DATA_TEMPR84[30] , 
        \R_DATA_TEMPR85[30] , \R_DATA_TEMPR86[30] , 
        \R_DATA_TEMPR87[30] , \R_DATA_TEMPR88[30] , 
        \R_DATA_TEMPR89[30] , \R_DATA_TEMPR90[30] , 
        \R_DATA_TEMPR91[30] , \R_DATA_TEMPR92[30] , 
        \R_DATA_TEMPR93[30] , \R_DATA_TEMPR94[30] , 
        \R_DATA_TEMPR95[30] , \R_DATA_TEMPR96[30] , 
        \R_DATA_TEMPR97[30] , \R_DATA_TEMPR98[30] , 
        \R_DATA_TEMPR99[30] , \R_DATA_TEMPR100[30] , 
        \R_DATA_TEMPR101[30] , \R_DATA_TEMPR102[30] , 
        \R_DATA_TEMPR103[30] , \R_DATA_TEMPR104[30] , 
        \R_DATA_TEMPR105[30] , \R_DATA_TEMPR106[30] , 
        \R_DATA_TEMPR107[30] , \R_DATA_TEMPR108[30] , 
        \R_DATA_TEMPR109[30] , \R_DATA_TEMPR110[30] , 
        \R_DATA_TEMPR111[30] , \R_DATA_TEMPR112[30] , 
        \R_DATA_TEMPR113[30] , \R_DATA_TEMPR114[30] , 
        \R_DATA_TEMPR115[30] , \R_DATA_TEMPR116[30] , 
        \R_DATA_TEMPR117[30] , \R_DATA_TEMPR118[30] , 
        \R_DATA_TEMPR119[30] , \R_DATA_TEMPR120[30] , 
        \R_DATA_TEMPR121[30] , \R_DATA_TEMPR122[30] , 
        \R_DATA_TEMPR123[30] , \R_DATA_TEMPR124[30] , 
        \R_DATA_TEMPR125[30] , \R_DATA_TEMPR126[30] , 
        \R_DATA_TEMPR127[30] , \R_DATA_TEMPR0[31] , 
        \R_DATA_TEMPR1[31] , \R_DATA_TEMPR2[31] , \R_DATA_TEMPR3[31] , 
        \R_DATA_TEMPR4[31] , \R_DATA_TEMPR5[31] , \R_DATA_TEMPR6[31] , 
        \R_DATA_TEMPR7[31] , \R_DATA_TEMPR8[31] , \R_DATA_TEMPR9[31] , 
        \R_DATA_TEMPR10[31] , \R_DATA_TEMPR11[31] , 
        \R_DATA_TEMPR12[31] , \R_DATA_TEMPR13[31] , 
        \R_DATA_TEMPR14[31] , \R_DATA_TEMPR15[31] , 
        \R_DATA_TEMPR16[31] , \R_DATA_TEMPR17[31] , 
        \R_DATA_TEMPR18[31] , \R_DATA_TEMPR19[31] , 
        \R_DATA_TEMPR20[31] , \R_DATA_TEMPR21[31] , 
        \R_DATA_TEMPR22[31] , \R_DATA_TEMPR23[31] , 
        \R_DATA_TEMPR24[31] , \R_DATA_TEMPR25[31] , 
        \R_DATA_TEMPR26[31] , \R_DATA_TEMPR27[31] , 
        \R_DATA_TEMPR28[31] , \R_DATA_TEMPR29[31] , 
        \R_DATA_TEMPR30[31] , \R_DATA_TEMPR31[31] , 
        \R_DATA_TEMPR32[31] , \R_DATA_TEMPR33[31] , 
        \R_DATA_TEMPR34[31] , \R_DATA_TEMPR35[31] , 
        \R_DATA_TEMPR36[31] , \R_DATA_TEMPR37[31] , 
        \R_DATA_TEMPR38[31] , \R_DATA_TEMPR39[31] , 
        \R_DATA_TEMPR40[31] , \R_DATA_TEMPR41[31] , 
        \R_DATA_TEMPR42[31] , \R_DATA_TEMPR43[31] , 
        \R_DATA_TEMPR44[31] , \R_DATA_TEMPR45[31] , 
        \R_DATA_TEMPR46[31] , \R_DATA_TEMPR47[31] , 
        \R_DATA_TEMPR48[31] , \R_DATA_TEMPR49[31] , 
        \R_DATA_TEMPR50[31] , \R_DATA_TEMPR51[31] , 
        \R_DATA_TEMPR52[31] , \R_DATA_TEMPR53[31] , 
        \R_DATA_TEMPR54[31] , \R_DATA_TEMPR55[31] , 
        \R_DATA_TEMPR56[31] , \R_DATA_TEMPR57[31] , 
        \R_DATA_TEMPR58[31] , \R_DATA_TEMPR59[31] , 
        \R_DATA_TEMPR60[31] , \R_DATA_TEMPR61[31] , 
        \R_DATA_TEMPR62[31] , \R_DATA_TEMPR63[31] , 
        \R_DATA_TEMPR64[31] , \R_DATA_TEMPR65[31] , 
        \R_DATA_TEMPR66[31] , \R_DATA_TEMPR67[31] , 
        \R_DATA_TEMPR68[31] , \R_DATA_TEMPR69[31] , 
        \R_DATA_TEMPR70[31] , \R_DATA_TEMPR71[31] , 
        \R_DATA_TEMPR72[31] , \R_DATA_TEMPR73[31] , 
        \R_DATA_TEMPR74[31] , \R_DATA_TEMPR75[31] , 
        \R_DATA_TEMPR76[31] , \R_DATA_TEMPR77[31] , 
        \R_DATA_TEMPR78[31] , \R_DATA_TEMPR79[31] , 
        \R_DATA_TEMPR80[31] , \R_DATA_TEMPR81[31] , 
        \R_DATA_TEMPR82[31] , \R_DATA_TEMPR83[31] , 
        \R_DATA_TEMPR84[31] , \R_DATA_TEMPR85[31] , 
        \R_DATA_TEMPR86[31] , \R_DATA_TEMPR87[31] , 
        \R_DATA_TEMPR88[31] , \R_DATA_TEMPR89[31] , 
        \R_DATA_TEMPR90[31] , \R_DATA_TEMPR91[31] , 
        \R_DATA_TEMPR92[31] , \R_DATA_TEMPR93[31] , 
        \R_DATA_TEMPR94[31] , \R_DATA_TEMPR95[31] , 
        \R_DATA_TEMPR96[31] , \R_DATA_TEMPR97[31] , 
        \R_DATA_TEMPR98[31] , \R_DATA_TEMPR99[31] , 
        \R_DATA_TEMPR100[31] , \R_DATA_TEMPR101[31] , 
        \R_DATA_TEMPR102[31] , \R_DATA_TEMPR103[31] , 
        \R_DATA_TEMPR104[31] , \R_DATA_TEMPR105[31] , 
        \R_DATA_TEMPR106[31] , \R_DATA_TEMPR107[31] , 
        \R_DATA_TEMPR108[31] , \R_DATA_TEMPR109[31] , 
        \R_DATA_TEMPR110[31] , \R_DATA_TEMPR111[31] , 
        \R_DATA_TEMPR112[31] , \R_DATA_TEMPR113[31] , 
        \R_DATA_TEMPR114[31] , \R_DATA_TEMPR115[31] , 
        \R_DATA_TEMPR116[31] , \R_DATA_TEMPR117[31] , 
        \R_DATA_TEMPR118[31] , \R_DATA_TEMPR119[31] , 
        \R_DATA_TEMPR120[31] , \R_DATA_TEMPR121[31] , 
        \R_DATA_TEMPR122[31] , \R_DATA_TEMPR123[31] , 
        \R_DATA_TEMPR124[31] , \R_DATA_TEMPR125[31] , 
        \R_DATA_TEMPR126[31] , \R_DATA_TEMPR127[31] , 
        \R_DATA_TEMPR0[32] , \R_DATA_TEMPR1[32] , \R_DATA_TEMPR2[32] , 
        \R_DATA_TEMPR3[32] , \R_DATA_TEMPR4[32] , \R_DATA_TEMPR5[32] , 
        \R_DATA_TEMPR6[32] , \R_DATA_TEMPR7[32] , \R_DATA_TEMPR8[32] , 
        \R_DATA_TEMPR9[32] , \R_DATA_TEMPR10[32] , 
        \R_DATA_TEMPR11[32] , \R_DATA_TEMPR12[32] , 
        \R_DATA_TEMPR13[32] , \R_DATA_TEMPR14[32] , 
        \R_DATA_TEMPR15[32] , \R_DATA_TEMPR16[32] , 
        \R_DATA_TEMPR17[32] , \R_DATA_TEMPR18[32] , 
        \R_DATA_TEMPR19[32] , \R_DATA_TEMPR20[32] , 
        \R_DATA_TEMPR21[32] , \R_DATA_TEMPR22[32] , 
        \R_DATA_TEMPR23[32] , \R_DATA_TEMPR24[32] , 
        \R_DATA_TEMPR25[32] , \R_DATA_TEMPR26[32] , 
        \R_DATA_TEMPR27[32] , \R_DATA_TEMPR28[32] , 
        \R_DATA_TEMPR29[32] , \R_DATA_TEMPR30[32] , 
        \R_DATA_TEMPR31[32] , \R_DATA_TEMPR32[32] , 
        \R_DATA_TEMPR33[32] , \R_DATA_TEMPR34[32] , 
        \R_DATA_TEMPR35[32] , \R_DATA_TEMPR36[32] , 
        \R_DATA_TEMPR37[32] , \R_DATA_TEMPR38[32] , 
        \R_DATA_TEMPR39[32] , \R_DATA_TEMPR40[32] , 
        \R_DATA_TEMPR41[32] , \R_DATA_TEMPR42[32] , 
        \R_DATA_TEMPR43[32] , \R_DATA_TEMPR44[32] , 
        \R_DATA_TEMPR45[32] , \R_DATA_TEMPR46[32] , 
        \R_DATA_TEMPR47[32] , \R_DATA_TEMPR48[32] , 
        \R_DATA_TEMPR49[32] , \R_DATA_TEMPR50[32] , 
        \R_DATA_TEMPR51[32] , \R_DATA_TEMPR52[32] , 
        \R_DATA_TEMPR53[32] , \R_DATA_TEMPR54[32] , 
        \R_DATA_TEMPR55[32] , \R_DATA_TEMPR56[32] , 
        \R_DATA_TEMPR57[32] , \R_DATA_TEMPR58[32] , 
        \R_DATA_TEMPR59[32] , \R_DATA_TEMPR60[32] , 
        \R_DATA_TEMPR61[32] , \R_DATA_TEMPR62[32] , 
        \R_DATA_TEMPR63[32] , \R_DATA_TEMPR64[32] , 
        \R_DATA_TEMPR65[32] , \R_DATA_TEMPR66[32] , 
        \R_DATA_TEMPR67[32] , \R_DATA_TEMPR68[32] , 
        \R_DATA_TEMPR69[32] , \R_DATA_TEMPR70[32] , 
        \R_DATA_TEMPR71[32] , \R_DATA_TEMPR72[32] , 
        \R_DATA_TEMPR73[32] , \R_DATA_TEMPR74[32] , 
        \R_DATA_TEMPR75[32] , \R_DATA_TEMPR76[32] , 
        \R_DATA_TEMPR77[32] , \R_DATA_TEMPR78[32] , 
        \R_DATA_TEMPR79[32] , \R_DATA_TEMPR80[32] , 
        \R_DATA_TEMPR81[32] , \R_DATA_TEMPR82[32] , 
        \R_DATA_TEMPR83[32] , \R_DATA_TEMPR84[32] , 
        \R_DATA_TEMPR85[32] , \R_DATA_TEMPR86[32] , 
        \R_DATA_TEMPR87[32] , \R_DATA_TEMPR88[32] , 
        \R_DATA_TEMPR89[32] , \R_DATA_TEMPR90[32] , 
        \R_DATA_TEMPR91[32] , \R_DATA_TEMPR92[32] , 
        \R_DATA_TEMPR93[32] , \R_DATA_TEMPR94[32] , 
        \R_DATA_TEMPR95[32] , \R_DATA_TEMPR96[32] , 
        \R_DATA_TEMPR97[32] , \R_DATA_TEMPR98[32] , 
        \R_DATA_TEMPR99[32] , \R_DATA_TEMPR100[32] , 
        \R_DATA_TEMPR101[32] , \R_DATA_TEMPR102[32] , 
        \R_DATA_TEMPR103[32] , \R_DATA_TEMPR104[32] , 
        \R_DATA_TEMPR105[32] , \R_DATA_TEMPR106[32] , 
        \R_DATA_TEMPR107[32] , \R_DATA_TEMPR108[32] , 
        \R_DATA_TEMPR109[32] , \R_DATA_TEMPR110[32] , 
        \R_DATA_TEMPR111[32] , \R_DATA_TEMPR112[32] , 
        \R_DATA_TEMPR113[32] , \R_DATA_TEMPR114[32] , 
        \R_DATA_TEMPR115[32] , \R_DATA_TEMPR116[32] , 
        \R_DATA_TEMPR117[32] , \R_DATA_TEMPR118[32] , 
        \R_DATA_TEMPR119[32] , \R_DATA_TEMPR120[32] , 
        \R_DATA_TEMPR121[32] , \R_DATA_TEMPR122[32] , 
        \R_DATA_TEMPR123[32] , \R_DATA_TEMPR124[32] , 
        \R_DATA_TEMPR125[32] , \R_DATA_TEMPR126[32] , 
        \R_DATA_TEMPR127[32] , \R_DATA_TEMPR0[33] , 
        \R_DATA_TEMPR1[33] , \R_DATA_TEMPR2[33] , \R_DATA_TEMPR3[33] , 
        \R_DATA_TEMPR4[33] , \R_DATA_TEMPR5[33] , \R_DATA_TEMPR6[33] , 
        \R_DATA_TEMPR7[33] , \R_DATA_TEMPR8[33] , \R_DATA_TEMPR9[33] , 
        \R_DATA_TEMPR10[33] , \R_DATA_TEMPR11[33] , 
        \R_DATA_TEMPR12[33] , \R_DATA_TEMPR13[33] , 
        \R_DATA_TEMPR14[33] , \R_DATA_TEMPR15[33] , 
        \R_DATA_TEMPR16[33] , \R_DATA_TEMPR17[33] , 
        \R_DATA_TEMPR18[33] , \R_DATA_TEMPR19[33] , 
        \R_DATA_TEMPR20[33] , \R_DATA_TEMPR21[33] , 
        \R_DATA_TEMPR22[33] , \R_DATA_TEMPR23[33] , 
        \R_DATA_TEMPR24[33] , \R_DATA_TEMPR25[33] , 
        \R_DATA_TEMPR26[33] , \R_DATA_TEMPR27[33] , 
        \R_DATA_TEMPR28[33] , \R_DATA_TEMPR29[33] , 
        \R_DATA_TEMPR30[33] , \R_DATA_TEMPR31[33] , 
        \R_DATA_TEMPR32[33] , \R_DATA_TEMPR33[33] , 
        \R_DATA_TEMPR34[33] , \R_DATA_TEMPR35[33] , 
        \R_DATA_TEMPR36[33] , \R_DATA_TEMPR37[33] , 
        \R_DATA_TEMPR38[33] , \R_DATA_TEMPR39[33] , 
        \R_DATA_TEMPR40[33] , \R_DATA_TEMPR41[33] , 
        \R_DATA_TEMPR42[33] , \R_DATA_TEMPR43[33] , 
        \R_DATA_TEMPR44[33] , \R_DATA_TEMPR45[33] , 
        \R_DATA_TEMPR46[33] , \R_DATA_TEMPR47[33] , 
        \R_DATA_TEMPR48[33] , \R_DATA_TEMPR49[33] , 
        \R_DATA_TEMPR50[33] , \R_DATA_TEMPR51[33] , 
        \R_DATA_TEMPR52[33] , \R_DATA_TEMPR53[33] , 
        \R_DATA_TEMPR54[33] , \R_DATA_TEMPR55[33] , 
        \R_DATA_TEMPR56[33] , \R_DATA_TEMPR57[33] , 
        \R_DATA_TEMPR58[33] , \R_DATA_TEMPR59[33] , 
        \R_DATA_TEMPR60[33] , \R_DATA_TEMPR61[33] , 
        \R_DATA_TEMPR62[33] , \R_DATA_TEMPR63[33] , 
        \R_DATA_TEMPR64[33] , \R_DATA_TEMPR65[33] , 
        \R_DATA_TEMPR66[33] , \R_DATA_TEMPR67[33] , 
        \R_DATA_TEMPR68[33] , \R_DATA_TEMPR69[33] , 
        \R_DATA_TEMPR70[33] , \R_DATA_TEMPR71[33] , 
        \R_DATA_TEMPR72[33] , \R_DATA_TEMPR73[33] , 
        \R_DATA_TEMPR74[33] , \R_DATA_TEMPR75[33] , 
        \R_DATA_TEMPR76[33] , \R_DATA_TEMPR77[33] , 
        \R_DATA_TEMPR78[33] , \R_DATA_TEMPR79[33] , 
        \R_DATA_TEMPR80[33] , \R_DATA_TEMPR81[33] , 
        \R_DATA_TEMPR82[33] , \R_DATA_TEMPR83[33] , 
        \R_DATA_TEMPR84[33] , \R_DATA_TEMPR85[33] , 
        \R_DATA_TEMPR86[33] , \R_DATA_TEMPR87[33] , 
        \R_DATA_TEMPR88[33] , \R_DATA_TEMPR89[33] , 
        \R_DATA_TEMPR90[33] , \R_DATA_TEMPR91[33] , 
        \R_DATA_TEMPR92[33] , \R_DATA_TEMPR93[33] , 
        \R_DATA_TEMPR94[33] , \R_DATA_TEMPR95[33] , 
        \R_DATA_TEMPR96[33] , \R_DATA_TEMPR97[33] , 
        \R_DATA_TEMPR98[33] , \R_DATA_TEMPR99[33] , 
        \R_DATA_TEMPR100[33] , \R_DATA_TEMPR101[33] , 
        \R_DATA_TEMPR102[33] , \R_DATA_TEMPR103[33] , 
        \R_DATA_TEMPR104[33] , \R_DATA_TEMPR105[33] , 
        \R_DATA_TEMPR106[33] , \R_DATA_TEMPR107[33] , 
        \R_DATA_TEMPR108[33] , \R_DATA_TEMPR109[33] , 
        \R_DATA_TEMPR110[33] , \R_DATA_TEMPR111[33] , 
        \R_DATA_TEMPR112[33] , \R_DATA_TEMPR113[33] , 
        \R_DATA_TEMPR114[33] , \R_DATA_TEMPR115[33] , 
        \R_DATA_TEMPR116[33] , \R_DATA_TEMPR117[33] , 
        \R_DATA_TEMPR118[33] , \R_DATA_TEMPR119[33] , 
        \R_DATA_TEMPR120[33] , \R_DATA_TEMPR121[33] , 
        \R_DATA_TEMPR122[33] , \R_DATA_TEMPR123[33] , 
        \R_DATA_TEMPR124[33] , \R_DATA_TEMPR125[33] , 
        \R_DATA_TEMPR126[33] , \R_DATA_TEMPR127[33] , 
        \R_DATA_TEMPR0[34] , \R_DATA_TEMPR1[34] , \R_DATA_TEMPR2[34] , 
        \R_DATA_TEMPR3[34] , \R_DATA_TEMPR4[34] , \R_DATA_TEMPR5[34] , 
        \R_DATA_TEMPR6[34] , \R_DATA_TEMPR7[34] , \R_DATA_TEMPR8[34] , 
        \R_DATA_TEMPR9[34] , \R_DATA_TEMPR10[34] , 
        \R_DATA_TEMPR11[34] , \R_DATA_TEMPR12[34] , 
        \R_DATA_TEMPR13[34] , \R_DATA_TEMPR14[34] , 
        \R_DATA_TEMPR15[34] , \R_DATA_TEMPR16[34] , 
        \R_DATA_TEMPR17[34] , \R_DATA_TEMPR18[34] , 
        \R_DATA_TEMPR19[34] , \R_DATA_TEMPR20[34] , 
        \R_DATA_TEMPR21[34] , \R_DATA_TEMPR22[34] , 
        \R_DATA_TEMPR23[34] , \R_DATA_TEMPR24[34] , 
        \R_DATA_TEMPR25[34] , \R_DATA_TEMPR26[34] , 
        \R_DATA_TEMPR27[34] , \R_DATA_TEMPR28[34] , 
        \R_DATA_TEMPR29[34] , \R_DATA_TEMPR30[34] , 
        \R_DATA_TEMPR31[34] , \R_DATA_TEMPR32[34] , 
        \R_DATA_TEMPR33[34] , \R_DATA_TEMPR34[34] , 
        \R_DATA_TEMPR35[34] , \R_DATA_TEMPR36[34] , 
        \R_DATA_TEMPR37[34] , \R_DATA_TEMPR38[34] , 
        \R_DATA_TEMPR39[34] , \R_DATA_TEMPR40[34] , 
        \R_DATA_TEMPR41[34] , \R_DATA_TEMPR42[34] , 
        \R_DATA_TEMPR43[34] , \R_DATA_TEMPR44[34] , 
        \R_DATA_TEMPR45[34] , \R_DATA_TEMPR46[34] , 
        \R_DATA_TEMPR47[34] , \R_DATA_TEMPR48[34] , 
        \R_DATA_TEMPR49[34] , \R_DATA_TEMPR50[34] , 
        \R_DATA_TEMPR51[34] , \R_DATA_TEMPR52[34] , 
        \R_DATA_TEMPR53[34] , \R_DATA_TEMPR54[34] , 
        \R_DATA_TEMPR55[34] , \R_DATA_TEMPR56[34] , 
        \R_DATA_TEMPR57[34] , \R_DATA_TEMPR58[34] , 
        \R_DATA_TEMPR59[34] , \R_DATA_TEMPR60[34] , 
        \R_DATA_TEMPR61[34] , \R_DATA_TEMPR62[34] , 
        \R_DATA_TEMPR63[34] , \R_DATA_TEMPR64[34] , 
        \R_DATA_TEMPR65[34] , \R_DATA_TEMPR66[34] , 
        \R_DATA_TEMPR67[34] , \R_DATA_TEMPR68[34] , 
        \R_DATA_TEMPR69[34] , \R_DATA_TEMPR70[34] , 
        \R_DATA_TEMPR71[34] , \R_DATA_TEMPR72[34] , 
        \R_DATA_TEMPR73[34] , \R_DATA_TEMPR74[34] , 
        \R_DATA_TEMPR75[34] , \R_DATA_TEMPR76[34] , 
        \R_DATA_TEMPR77[34] , \R_DATA_TEMPR78[34] , 
        \R_DATA_TEMPR79[34] , \R_DATA_TEMPR80[34] , 
        \R_DATA_TEMPR81[34] , \R_DATA_TEMPR82[34] , 
        \R_DATA_TEMPR83[34] , \R_DATA_TEMPR84[34] , 
        \R_DATA_TEMPR85[34] , \R_DATA_TEMPR86[34] , 
        \R_DATA_TEMPR87[34] , \R_DATA_TEMPR88[34] , 
        \R_DATA_TEMPR89[34] , \R_DATA_TEMPR90[34] , 
        \R_DATA_TEMPR91[34] , \R_DATA_TEMPR92[34] , 
        \R_DATA_TEMPR93[34] , \R_DATA_TEMPR94[34] , 
        \R_DATA_TEMPR95[34] , \R_DATA_TEMPR96[34] , 
        \R_DATA_TEMPR97[34] , \R_DATA_TEMPR98[34] , 
        \R_DATA_TEMPR99[34] , \R_DATA_TEMPR100[34] , 
        \R_DATA_TEMPR101[34] , \R_DATA_TEMPR102[34] , 
        \R_DATA_TEMPR103[34] , \R_DATA_TEMPR104[34] , 
        \R_DATA_TEMPR105[34] , \R_DATA_TEMPR106[34] , 
        \R_DATA_TEMPR107[34] , \R_DATA_TEMPR108[34] , 
        \R_DATA_TEMPR109[34] , \R_DATA_TEMPR110[34] , 
        \R_DATA_TEMPR111[34] , \R_DATA_TEMPR112[34] , 
        \R_DATA_TEMPR113[34] , \R_DATA_TEMPR114[34] , 
        \R_DATA_TEMPR115[34] , \R_DATA_TEMPR116[34] , 
        \R_DATA_TEMPR117[34] , \R_DATA_TEMPR118[34] , 
        \R_DATA_TEMPR119[34] , \R_DATA_TEMPR120[34] , 
        \R_DATA_TEMPR121[34] , \R_DATA_TEMPR122[34] , 
        \R_DATA_TEMPR123[34] , \R_DATA_TEMPR124[34] , 
        \R_DATA_TEMPR125[34] , \R_DATA_TEMPR126[34] , 
        \R_DATA_TEMPR127[34] , \R_DATA_TEMPR0[35] , 
        \R_DATA_TEMPR1[35] , \R_DATA_TEMPR2[35] , \R_DATA_TEMPR3[35] , 
        \R_DATA_TEMPR4[35] , \R_DATA_TEMPR5[35] , \R_DATA_TEMPR6[35] , 
        \R_DATA_TEMPR7[35] , \R_DATA_TEMPR8[35] , \R_DATA_TEMPR9[35] , 
        \R_DATA_TEMPR10[35] , \R_DATA_TEMPR11[35] , 
        \R_DATA_TEMPR12[35] , \R_DATA_TEMPR13[35] , 
        \R_DATA_TEMPR14[35] , \R_DATA_TEMPR15[35] , 
        \R_DATA_TEMPR16[35] , \R_DATA_TEMPR17[35] , 
        \R_DATA_TEMPR18[35] , \R_DATA_TEMPR19[35] , 
        \R_DATA_TEMPR20[35] , \R_DATA_TEMPR21[35] , 
        \R_DATA_TEMPR22[35] , \R_DATA_TEMPR23[35] , 
        \R_DATA_TEMPR24[35] , \R_DATA_TEMPR25[35] , 
        \R_DATA_TEMPR26[35] , \R_DATA_TEMPR27[35] , 
        \R_DATA_TEMPR28[35] , \R_DATA_TEMPR29[35] , 
        \R_DATA_TEMPR30[35] , \R_DATA_TEMPR31[35] , 
        \R_DATA_TEMPR32[35] , \R_DATA_TEMPR33[35] , 
        \R_DATA_TEMPR34[35] , \R_DATA_TEMPR35[35] , 
        \R_DATA_TEMPR36[35] , \R_DATA_TEMPR37[35] , 
        \R_DATA_TEMPR38[35] , \R_DATA_TEMPR39[35] , 
        \R_DATA_TEMPR40[35] , \R_DATA_TEMPR41[35] , 
        \R_DATA_TEMPR42[35] , \R_DATA_TEMPR43[35] , 
        \R_DATA_TEMPR44[35] , \R_DATA_TEMPR45[35] , 
        \R_DATA_TEMPR46[35] , \R_DATA_TEMPR47[35] , 
        \R_DATA_TEMPR48[35] , \R_DATA_TEMPR49[35] , 
        \R_DATA_TEMPR50[35] , \R_DATA_TEMPR51[35] , 
        \R_DATA_TEMPR52[35] , \R_DATA_TEMPR53[35] , 
        \R_DATA_TEMPR54[35] , \R_DATA_TEMPR55[35] , 
        \R_DATA_TEMPR56[35] , \R_DATA_TEMPR57[35] , 
        \R_DATA_TEMPR58[35] , \R_DATA_TEMPR59[35] , 
        \R_DATA_TEMPR60[35] , \R_DATA_TEMPR61[35] , 
        \R_DATA_TEMPR62[35] , \R_DATA_TEMPR63[35] , 
        \R_DATA_TEMPR64[35] , \R_DATA_TEMPR65[35] , 
        \R_DATA_TEMPR66[35] , \R_DATA_TEMPR67[35] , 
        \R_DATA_TEMPR68[35] , \R_DATA_TEMPR69[35] , 
        \R_DATA_TEMPR70[35] , \R_DATA_TEMPR71[35] , 
        \R_DATA_TEMPR72[35] , \R_DATA_TEMPR73[35] , 
        \R_DATA_TEMPR74[35] , \R_DATA_TEMPR75[35] , 
        \R_DATA_TEMPR76[35] , \R_DATA_TEMPR77[35] , 
        \R_DATA_TEMPR78[35] , \R_DATA_TEMPR79[35] , 
        \R_DATA_TEMPR80[35] , \R_DATA_TEMPR81[35] , 
        \R_DATA_TEMPR82[35] , \R_DATA_TEMPR83[35] , 
        \R_DATA_TEMPR84[35] , \R_DATA_TEMPR85[35] , 
        \R_DATA_TEMPR86[35] , \R_DATA_TEMPR87[35] , 
        \R_DATA_TEMPR88[35] , \R_DATA_TEMPR89[35] , 
        \R_DATA_TEMPR90[35] , \R_DATA_TEMPR91[35] , 
        \R_DATA_TEMPR92[35] , \R_DATA_TEMPR93[35] , 
        \R_DATA_TEMPR94[35] , \R_DATA_TEMPR95[35] , 
        \R_DATA_TEMPR96[35] , \R_DATA_TEMPR97[35] , 
        \R_DATA_TEMPR98[35] , \R_DATA_TEMPR99[35] , 
        \R_DATA_TEMPR100[35] , \R_DATA_TEMPR101[35] , 
        \R_DATA_TEMPR102[35] , \R_DATA_TEMPR103[35] , 
        \R_DATA_TEMPR104[35] , \R_DATA_TEMPR105[35] , 
        \R_DATA_TEMPR106[35] , \R_DATA_TEMPR107[35] , 
        \R_DATA_TEMPR108[35] , \R_DATA_TEMPR109[35] , 
        \R_DATA_TEMPR110[35] , \R_DATA_TEMPR111[35] , 
        \R_DATA_TEMPR112[35] , \R_DATA_TEMPR113[35] , 
        \R_DATA_TEMPR114[35] , \R_DATA_TEMPR115[35] , 
        \R_DATA_TEMPR116[35] , \R_DATA_TEMPR117[35] , 
        \R_DATA_TEMPR118[35] , \R_DATA_TEMPR119[35] , 
        \R_DATA_TEMPR120[35] , \R_DATA_TEMPR121[35] , 
        \R_DATA_TEMPR122[35] , \R_DATA_TEMPR123[35] , 
        \R_DATA_TEMPR124[35] , \R_DATA_TEMPR125[35] , 
        \R_DATA_TEMPR126[35] , \R_DATA_TEMPR127[35] , 
        \R_DATA_TEMPR0[36] , \R_DATA_TEMPR1[36] , \R_DATA_TEMPR2[36] , 
        \R_DATA_TEMPR3[36] , \R_DATA_TEMPR4[36] , \R_DATA_TEMPR5[36] , 
        \R_DATA_TEMPR6[36] , \R_DATA_TEMPR7[36] , \R_DATA_TEMPR8[36] , 
        \R_DATA_TEMPR9[36] , \R_DATA_TEMPR10[36] , 
        \R_DATA_TEMPR11[36] , \R_DATA_TEMPR12[36] , 
        \R_DATA_TEMPR13[36] , \R_DATA_TEMPR14[36] , 
        \R_DATA_TEMPR15[36] , \R_DATA_TEMPR16[36] , 
        \R_DATA_TEMPR17[36] , \R_DATA_TEMPR18[36] , 
        \R_DATA_TEMPR19[36] , \R_DATA_TEMPR20[36] , 
        \R_DATA_TEMPR21[36] , \R_DATA_TEMPR22[36] , 
        \R_DATA_TEMPR23[36] , \R_DATA_TEMPR24[36] , 
        \R_DATA_TEMPR25[36] , \R_DATA_TEMPR26[36] , 
        \R_DATA_TEMPR27[36] , \R_DATA_TEMPR28[36] , 
        \R_DATA_TEMPR29[36] , \R_DATA_TEMPR30[36] , 
        \R_DATA_TEMPR31[36] , \R_DATA_TEMPR32[36] , 
        \R_DATA_TEMPR33[36] , \R_DATA_TEMPR34[36] , 
        \R_DATA_TEMPR35[36] , \R_DATA_TEMPR36[36] , 
        \R_DATA_TEMPR37[36] , \R_DATA_TEMPR38[36] , 
        \R_DATA_TEMPR39[36] , \R_DATA_TEMPR40[36] , 
        \R_DATA_TEMPR41[36] , \R_DATA_TEMPR42[36] , 
        \R_DATA_TEMPR43[36] , \R_DATA_TEMPR44[36] , 
        \R_DATA_TEMPR45[36] , \R_DATA_TEMPR46[36] , 
        \R_DATA_TEMPR47[36] , \R_DATA_TEMPR48[36] , 
        \R_DATA_TEMPR49[36] , \R_DATA_TEMPR50[36] , 
        \R_DATA_TEMPR51[36] , \R_DATA_TEMPR52[36] , 
        \R_DATA_TEMPR53[36] , \R_DATA_TEMPR54[36] , 
        \R_DATA_TEMPR55[36] , \R_DATA_TEMPR56[36] , 
        \R_DATA_TEMPR57[36] , \R_DATA_TEMPR58[36] , 
        \R_DATA_TEMPR59[36] , \R_DATA_TEMPR60[36] , 
        \R_DATA_TEMPR61[36] , \R_DATA_TEMPR62[36] , 
        \R_DATA_TEMPR63[36] , \R_DATA_TEMPR64[36] , 
        \R_DATA_TEMPR65[36] , \R_DATA_TEMPR66[36] , 
        \R_DATA_TEMPR67[36] , \R_DATA_TEMPR68[36] , 
        \R_DATA_TEMPR69[36] , \R_DATA_TEMPR70[36] , 
        \R_DATA_TEMPR71[36] , \R_DATA_TEMPR72[36] , 
        \R_DATA_TEMPR73[36] , \R_DATA_TEMPR74[36] , 
        \R_DATA_TEMPR75[36] , \R_DATA_TEMPR76[36] , 
        \R_DATA_TEMPR77[36] , \R_DATA_TEMPR78[36] , 
        \R_DATA_TEMPR79[36] , \R_DATA_TEMPR80[36] , 
        \R_DATA_TEMPR81[36] , \R_DATA_TEMPR82[36] , 
        \R_DATA_TEMPR83[36] , \R_DATA_TEMPR84[36] , 
        \R_DATA_TEMPR85[36] , \R_DATA_TEMPR86[36] , 
        \R_DATA_TEMPR87[36] , \R_DATA_TEMPR88[36] , 
        \R_DATA_TEMPR89[36] , \R_DATA_TEMPR90[36] , 
        \R_DATA_TEMPR91[36] , \R_DATA_TEMPR92[36] , 
        \R_DATA_TEMPR93[36] , \R_DATA_TEMPR94[36] , 
        \R_DATA_TEMPR95[36] , \R_DATA_TEMPR96[36] , 
        \R_DATA_TEMPR97[36] , \R_DATA_TEMPR98[36] , 
        \R_DATA_TEMPR99[36] , \R_DATA_TEMPR100[36] , 
        \R_DATA_TEMPR101[36] , \R_DATA_TEMPR102[36] , 
        \R_DATA_TEMPR103[36] , \R_DATA_TEMPR104[36] , 
        \R_DATA_TEMPR105[36] , \R_DATA_TEMPR106[36] , 
        \R_DATA_TEMPR107[36] , \R_DATA_TEMPR108[36] , 
        \R_DATA_TEMPR109[36] , \R_DATA_TEMPR110[36] , 
        \R_DATA_TEMPR111[36] , \R_DATA_TEMPR112[36] , 
        \R_DATA_TEMPR113[36] , \R_DATA_TEMPR114[36] , 
        \R_DATA_TEMPR115[36] , \R_DATA_TEMPR116[36] , 
        \R_DATA_TEMPR117[36] , \R_DATA_TEMPR118[36] , 
        \R_DATA_TEMPR119[36] , \R_DATA_TEMPR120[36] , 
        \R_DATA_TEMPR121[36] , \R_DATA_TEMPR122[36] , 
        \R_DATA_TEMPR123[36] , \R_DATA_TEMPR124[36] , 
        \R_DATA_TEMPR125[36] , \R_DATA_TEMPR126[36] , 
        \R_DATA_TEMPR127[36] , \R_DATA_TEMPR0[37] , 
        \R_DATA_TEMPR1[37] , \R_DATA_TEMPR2[37] , \R_DATA_TEMPR3[37] , 
        \R_DATA_TEMPR4[37] , \R_DATA_TEMPR5[37] , \R_DATA_TEMPR6[37] , 
        \R_DATA_TEMPR7[37] , \R_DATA_TEMPR8[37] , \R_DATA_TEMPR9[37] , 
        \R_DATA_TEMPR10[37] , \R_DATA_TEMPR11[37] , 
        \R_DATA_TEMPR12[37] , \R_DATA_TEMPR13[37] , 
        \R_DATA_TEMPR14[37] , \R_DATA_TEMPR15[37] , 
        \R_DATA_TEMPR16[37] , \R_DATA_TEMPR17[37] , 
        \R_DATA_TEMPR18[37] , \R_DATA_TEMPR19[37] , 
        \R_DATA_TEMPR20[37] , \R_DATA_TEMPR21[37] , 
        \R_DATA_TEMPR22[37] , \R_DATA_TEMPR23[37] , 
        \R_DATA_TEMPR24[37] , \R_DATA_TEMPR25[37] , 
        \R_DATA_TEMPR26[37] , \R_DATA_TEMPR27[37] , 
        \R_DATA_TEMPR28[37] , \R_DATA_TEMPR29[37] , 
        \R_DATA_TEMPR30[37] , \R_DATA_TEMPR31[37] , 
        \R_DATA_TEMPR32[37] , \R_DATA_TEMPR33[37] , 
        \R_DATA_TEMPR34[37] , \R_DATA_TEMPR35[37] , 
        \R_DATA_TEMPR36[37] , \R_DATA_TEMPR37[37] , 
        \R_DATA_TEMPR38[37] , \R_DATA_TEMPR39[37] , 
        \R_DATA_TEMPR40[37] , \R_DATA_TEMPR41[37] , 
        \R_DATA_TEMPR42[37] , \R_DATA_TEMPR43[37] , 
        \R_DATA_TEMPR44[37] , \R_DATA_TEMPR45[37] , 
        \R_DATA_TEMPR46[37] , \R_DATA_TEMPR47[37] , 
        \R_DATA_TEMPR48[37] , \R_DATA_TEMPR49[37] , 
        \R_DATA_TEMPR50[37] , \R_DATA_TEMPR51[37] , 
        \R_DATA_TEMPR52[37] , \R_DATA_TEMPR53[37] , 
        \R_DATA_TEMPR54[37] , \R_DATA_TEMPR55[37] , 
        \R_DATA_TEMPR56[37] , \R_DATA_TEMPR57[37] , 
        \R_DATA_TEMPR58[37] , \R_DATA_TEMPR59[37] , 
        \R_DATA_TEMPR60[37] , \R_DATA_TEMPR61[37] , 
        \R_DATA_TEMPR62[37] , \R_DATA_TEMPR63[37] , 
        \R_DATA_TEMPR64[37] , \R_DATA_TEMPR65[37] , 
        \R_DATA_TEMPR66[37] , \R_DATA_TEMPR67[37] , 
        \R_DATA_TEMPR68[37] , \R_DATA_TEMPR69[37] , 
        \R_DATA_TEMPR70[37] , \R_DATA_TEMPR71[37] , 
        \R_DATA_TEMPR72[37] , \R_DATA_TEMPR73[37] , 
        \R_DATA_TEMPR74[37] , \R_DATA_TEMPR75[37] , 
        \R_DATA_TEMPR76[37] , \R_DATA_TEMPR77[37] , 
        \R_DATA_TEMPR78[37] , \R_DATA_TEMPR79[37] , 
        \R_DATA_TEMPR80[37] , \R_DATA_TEMPR81[37] , 
        \R_DATA_TEMPR82[37] , \R_DATA_TEMPR83[37] , 
        \R_DATA_TEMPR84[37] , \R_DATA_TEMPR85[37] , 
        \R_DATA_TEMPR86[37] , \R_DATA_TEMPR87[37] , 
        \R_DATA_TEMPR88[37] , \R_DATA_TEMPR89[37] , 
        \R_DATA_TEMPR90[37] , \R_DATA_TEMPR91[37] , 
        \R_DATA_TEMPR92[37] , \R_DATA_TEMPR93[37] , 
        \R_DATA_TEMPR94[37] , \R_DATA_TEMPR95[37] , 
        \R_DATA_TEMPR96[37] , \R_DATA_TEMPR97[37] , 
        \R_DATA_TEMPR98[37] , \R_DATA_TEMPR99[37] , 
        \R_DATA_TEMPR100[37] , \R_DATA_TEMPR101[37] , 
        \R_DATA_TEMPR102[37] , \R_DATA_TEMPR103[37] , 
        \R_DATA_TEMPR104[37] , \R_DATA_TEMPR105[37] , 
        \R_DATA_TEMPR106[37] , \R_DATA_TEMPR107[37] , 
        \R_DATA_TEMPR108[37] , \R_DATA_TEMPR109[37] , 
        \R_DATA_TEMPR110[37] , \R_DATA_TEMPR111[37] , 
        \R_DATA_TEMPR112[37] , \R_DATA_TEMPR113[37] , 
        \R_DATA_TEMPR114[37] , \R_DATA_TEMPR115[37] , 
        \R_DATA_TEMPR116[37] , \R_DATA_TEMPR117[37] , 
        \R_DATA_TEMPR118[37] , \R_DATA_TEMPR119[37] , 
        \R_DATA_TEMPR120[37] , \R_DATA_TEMPR121[37] , 
        \R_DATA_TEMPR122[37] , \R_DATA_TEMPR123[37] , 
        \R_DATA_TEMPR124[37] , \R_DATA_TEMPR125[37] , 
        \R_DATA_TEMPR126[37] , \R_DATA_TEMPR127[37] , 
        \R_DATA_TEMPR0[38] , \R_DATA_TEMPR1[38] , \R_DATA_TEMPR2[38] , 
        \R_DATA_TEMPR3[38] , \R_DATA_TEMPR4[38] , \R_DATA_TEMPR5[38] , 
        \R_DATA_TEMPR6[38] , \R_DATA_TEMPR7[38] , \R_DATA_TEMPR8[38] , 
        \R_DATA_TEMPR9[38] , \R_DATA_TEMPR10[38] , 
        \R_DATA_TEMPR11[38] , \R_DATA_TEMPR12[38] , 
        \R_DATA_TEMPR13[38] , \R_DATA_TEMPR14[38] , 
        \R_DATA_TEMPR15[38] , \R_DATA_TEMPR16[38] , 
        \R_DATA_TEMPR17[38] , \R_DATA_TEMPR18[38] , 
        \R_DATA_TEMPR19[38] , \R_DATA_TEMPR20[38] , 
        \R_DATA_TEMPR21[38] , \R_DATA_TEMPR22[38] , 
        \R_DATA_TEMPR23[38] , \R_DATA_TEMPR24[38] , 
        \R_DATA_TEMPR25[38] , \R_DATA_TEMPR26[38] , 
        \R_DATA_TEMPR27[38] , \R_DATA_TEMPR28[38] , 
        \R_DATA_TEMPR29[38] , \R_DATA_TEMPR30[38] , 
        \R_DATA_TEMPR31[38] , \R_DATA_TEMPR32[38] , 
        \R_DATA_TEMPR33[38] , \R_DATA_TEMPR34[38] , 
        \R_DATA_TEMPR35[38] , \R_DATA_TEMPR36[38] , 
        \R_DATA_TEMPR37[38] , \R_DATA_TEMPR38[38] , 
        \R_DATA_TEMPR39[38] , \R_DATA_TEMPR40[38] , 
        \R_DATA_TEMPR41[38] , \R_DATA_TEMPR42[38] , 
        \R_DATA_TEMPR43[38] , \R_DATA_TEMPR44[38] , 
        \R_DATA_TEMPR45[38] , \R_DATA_TEMPR46[38] , 
        \R_DATA_TEMPR47[38] , \R_DATA_TEMPR48[38] , 
        \R_DATA_TEMPR49[38] , \R_DATA_TEMPR50[38] , 
        \R_DATA_TEMPR51[38] , \R_DATA_TEMPR52[38] , 
        \R_DATA_TEMPR53[38] , \R_DATA_TEMPR54[38] , 
        \R_DATA_TEMPR55[38] , \R_DATA_TEMPR56[38] , 
        \R_DATA_TEMPR57[38] , \R_DATA_TEMPR58[38] , 
        \R_DATA_TEMPR59[38] , \R_DATA_TEMPR60[38] , 
        \R_DATA_TEMPR61[38] , \R_DATA_TEMPR62[38] , 
        \R_DATA_TEMPR63[38] , \R_DATA_TEMPR64[38] , 
        \R_DATA_TEMPR65[38] , \R_DATA_TEMPR66[38] , 
        \R_DATA_TEMPR67[38] , \R_DATA_TEMPR68[38] , 
        \R_DATA_TEMPR69[38] , \R_DATA_TEMPR70[38] , 
        \R_DATA_TEMPR71[38] , \R_DATA_TEMPR72[38] , 
        \R_DATA_TEMPR73[38] , \R_DATA_TEMPR74[38] , 
        \R_DATA_TEMPR75[38] , \R_DATA_TEMPR76[38] , 
        \R_DATA_TEMPR77[38] , \R_DATA_TEMPR78[38] , 
        \R_DATA_TEMPR79[38] , \R_DATA_TEMPR80[38] , 
        \R_DATA_TEMPR81[38] , \R_DATA_TEMPR82[38] , 
        \R_DATA_TEMPR83[38] , \R_DATA_TEMPR84[38] , 
        \R_DATA_TEMPR85[38] , \R_DATA_TEMPR86[38] , 
        \R_DATA_TEMPR87[38] , \R_DATA_TEMPR88[38] , 
        \R_DATA_TEMPR89[38] , \R_DATA_TEMPR90[38] , 
        \R_DATA_TEMPR91[38] , \R_DATA_TEMPR92[38] , 
        \R_DATA_TEMPR93[38] , \R_DATA_TEMPR94[38] , 
        \R_DATA_TEMPR95[38] , \R_DATA_TEMPR96[38] , 
        \R_DATA_TEMPR97[38] , \R_DATA_TEMPR98[38] , 
        \R_DATA_TEMPR99[38] , \R_DATA_TEMPR100[38] , 
        \R_DATA_TEMPR101[38] , \R_DATA_TEMPR102[38] , 
        \R_DATA_TEMPR103[38] , \R_DATA_TEMPR104[38] , 
        \R_DATA_TEMPR105[38] , \R_DATA_TEMPR106[38] , 
        \R_DATA_TEMPR107[38] , \R_DATA_TEMPR108[38] , 
        \R_DATA_TEMPR109[38] , \R_DATA_TEMPR110[38] , 
        \R_DATA_TEMPR111[38] , \R_DATA_TEMPR112[38] , 
        \R_DATA_TEMPR113[38] , \R_DATA_TEMPR114[38] , 
        \R_DATA_TEMPR115[38] , \R_DATA_TEMPR116[38] , 
        \R_DATA_TEMPR117[38] , \R_DATA_TEMPR118[38] , 
        \R_DATA_TEMPR119[38] , \R_DATA_TEMPR120[38] , 
        \R_DATA_TEMPR121[38] , \R_DATA_TEMPR122[38] , 
        \R_DATA_TEMPR123[38] , \R_DATA_TEMPR124[38] , 
        \R_DATA_TEMPR125[38] , \R_DATA_TEMPR126[38] , 
        \R_DATA_TEMPR127[38] , \R_DATA_TEMPR0[39] , 
        \R_DATA_TEMPR1[39] , \R_DATA_TEMPR2[39] , \R_DATA_TEMPR3[39] , 
        \R_DATA_TEMPR4[39] , \R_DATA_TEMPR5[39] , \R_DATA_TEMPR6[39] , 
        \R_DATA_TEMPR7[39] , \R_DATA_TEMPR8[39] , \R_DATA_TEMPR9[39] , 
        \R_DATA_TEMPR10[39] , \R_DATA_TEMPR11[39] , 
        \R_DATA_TEMPR12[39] , \R_DATA_TEMPR13[39] , 
        \R_DATA_TEMPR14[39] , \R_DATA_TEMPR15[39] , 
        \R_DATA_TEMPR16[39] , \R_DATA_TEMPR17[39] , 
        \R_DATA_TEMPR18[39] , \R_DATA_TEMPR19[39] , 
        \R_DATA_TEMPR20[39] , \R_DATA_TEMPR21[39] , 
        \R_DATA_TEMPR22[39] , \R_DATA_TEMPR23[39] , 
        \R_DATA_TEMPR24[39] , \R_DATA_TEMPR25[39] , 
        \R_DATA_TEMPR26[39] , \R_DATA_TEMPR27[39] , 
        \R_DATA_TEMPR28[39] , \R_DATA_TEMPR29[39] , 
        \R_DATA_TEMPR30[39] , \R_DATA_TEMPR31[39] , 
        \R_DATA_TEMPR32[39] , \R_DATA_TEMPR33[39] , 
        \R_DATA_TEMPR34[39] , \R_DATA_TEMPR35[39] , 
        \R_DATA_TEMPR36[39] , \R_DATA_TEMPR37[39] , 
        \R_DATA_TEMPR38[39] , \R_DATA_TEMPR39[39] , 
        \R_DATA_TEMPR40[39] , \R_DATA_TEMPR41[39] , 
        \R_DATA_TEMPR42[39] , \R_DATA_TEMPR43[39] , 
        \R_DATA_TEMPR44[39] , \R_DATA_TEMPR45[39] , 
        \R_DATA_TEMPR46[39] , \R_DATA_TEMPR47[39] , 
        \R_DATA_TEMPR48[39] , \R_DATA_TEMPR49[39] , 
        \R_DATA_TEMPR50[39] , \R_DATA_TEMPR51[39] , 
        \R_DATA_TEMPR52[39] , \R_DATA_TEMPR53[39] , 
        \R_DATA_TEMPR54[39] , \R_DATA_TEMPR55[39] , 
        \R_DATA_TEMPR56[39] , \R_DATA_TEMPR57[39] , 
        \R_DATA_TEMPR58[39] , \R_DATA_TEMPR59[39] , 
        \R_DATA_TEMPR60[39] , \R_DATA_TEMPR61[39] , 
        \R_DATA_TEMPR62[39] , \R_DATA_TEMPR63[39] , 
        \R_DATA_TEMPR64[39] , \R_DATA_TEMPR65[39] , 
        \R_DATA_TEMPR66[39] , \R_DATA_TEMPR67[39] , 
        \R_DATA_TEMPR68[39] , \R_DATA_TEMPR69[39] , 
        \R_DATA_TEMPR70[39] , \R_DATA_TEMPR71[39] , 
        \R_DATA_TEMPR72[39] , \R_DATA_TEMPR73[39] , 
        \R_DATA_TEMPR74[39] , \R_DATA_TEMPR75[39] , 
        \R_DATA_TEMPR76[39] , \R_DATA_TEMPR77[39] , 
        \R_DATA_TEMPR78[39] , \R_DATA_TEMPR79[39] , 
        \R_DATA_TEMPR80[39] , \R_DATA_TEMPR81[39] , 
        \R_DATA_TEMPR82[39] , \R_DATA_TEMPR83[39] , 
        \R_DATA_TEMPR84[39] , \R_DATA_TEMPR85[39] , 
        \R_DATA_TEMPR86[39] , \R_DATA_TEMPR87[39] , 
        \R_DATA_TEMPR88[39] , \R_DATA_TEMPR89[39] , 
        \R_DATA_TEMPR90[39] , \R_DATA_TEMPR91[39] , 
        \R_DATA_TEMPR92[39] , \R_DATA_TEMPR93[39] , 
        \R_DATA_TEMPR94[39] , \R_DATA_TEMPR95[39] , 
        \R_DATA_TEMPR96[39] , \R_DATA_TEMPR97[39] , 
        \R_DATA_TEMPR98[39] , \R_DATA_TEMPR99[39] , 
        \R_DATA_TEMPR100[39] , \R_DATA_TEMPR101[39] , 
        \R_DATA_TEMPR102[39] , \R_DATA_TEMPR103[39] , 
        \R_DATA_TEMPR104[39] , \R_DATA_TEMPR105[39] , 
        \R_DATA_TEMPR106[39] , \R_DATA_TEMPR107[39] , 
        \R_DATA_TEMPR108[39] , \R_DATA_TEMPR109[39] , 
        \R_DATA_TEMPR110[39] , \R_DATA_TEMPR111[39] , 
        \R_DATA_TEMPR112[39] , \R_DATA_TEMPR113[39] , 
        \R_DATA_TEMPR114[39] , \R_DATA_TEMPR115[39] , 
        \R_DATA_TEMPR116[39] , \R_DATA_TEMPR117[39] , 
        \R_DATA_TEMPR118[39] , \R_DATA_TEMPR119[39] , 
        \R_DATA_TEMPR120[39] , \R_DATA_TEMPR121[39] , 
        \R_DATA_TEMPR122[39] , \R_DATA_TEMPR123[39] , 
        \R_DATA_TEMPR124[39] , \R_DATA_TEMPR125[39] , 
        \R_DATA_TEMPR126[39] , \R_DATA_TEMPR127[39] , \BLKX0[0] , 
        \BLKY0[0] , \BLKX1[0] , \BLKY1[0] , \BLKX2[0] , \BLKX2[1] , 
        \BLKX2[2] , \BLKX2[3] , \BLKX2[4] , \BLKX2[5] , \BLKX2[6] , 
        \BLKX2[7] , \BLKX2[8] , \BLKX2[9] , \BLKX2[10] , \BLKX2[11] , 
        \BLKX2[12] , \BLKX2[13] , \BLKX2[14] , \BLKX2[15] , 
        \BLKX2[16] , \BLKX2[17] , \BLKX2[18] , \BLKX2[19] , 
        \BLKX2[20] , \BLKX2[21] , \BLKX2[22] , \BLKX2[23] , 
        \BLKX2[24] , \BLKX2[25] , \BLKX2[26] , \BLKX2[27] , 
        \BLKX2[28] , \BLKX2[29] , \BLKX2[30] , \BLKX2[31] , \BLKY2[0] , 
        \BLKY2[1] , \BLKY2[2] , \BLKY2[3] , \BLKY2[4] , \BLKY2[5] , 
        \BLKY2[6] , \BLKY2[7] , \BLKY2[8] , \BLKY2[9] , \BLKY2[10] , 
        \BLKY2[11] , \BLKY2[12] , \BLKY2[13] , \BLKY2[14] , 
        \BLKY2[15] , \BLKY2[16] , \BLKY2[17] , \BLKY2[18] , 
        \BLKY2[19] , \BLKY2[20] , \BLKY2[21] , \BLKY2[22] , 
        \BLKY2[23] , \BLKY2[24] , \BLKY2[25] , \BLKY2[26] , 
        \BLKY2[27] , \BLKY2[28] , \BLKY2[29] , \BLKY2[30] , 
        \BLKY2[31] , \ACCESS_BUSY[0][0] , \ACCESS_BUSY[1][0] , 
        \ACCESS_BUSY[2][0] , \ACCESS_BUSY[3][0] , \ACCESS_BUSY[4][0] , 
        \ACCESS_BUSY[5][0] , \ACCESS_BUSY[6][0] , \ACCESS_BUSY[7][0] , 
        \ACCESS_BUSY[8][0] , \ACCESS_BUSY[9][0] , \ACCESS_BUSY[10][0] , 
        \ACCESS_BUSY[11][0] , \ACCESS_BUSY[12][0] , 
        \ACCESS_BUSY[13][0] , \ACCESS_BUSY[14][0] , 
        \ACCESS_BUSY[15][0] , \ACCESS_BUSY[16][0] , 
        \ACCESS_BUSY[17][0] , \ACCESS_BUSY[18][0] , 
        \ACCESS_BUSY[19][0] , \ACCESS_BUSY[20][0] , 
        \ACCESS_BUSY[21][0] , \ACCESS_BUSY[22][0] , 
        \ACCESS_BUSY[23][0] , \ACCESS_BUSY[24][0] , 
        \ACCESS_BUSY[25][0] , \ACCESS_BUSY[26][0] , 
        \ACCESS_BUSY[27][0] , \ACCESS_BUSY[28][0] , 
        \ACCESS_BUSY[29][0] , \ACCESS_BUSY[30][0] , 
        \ACCESS_BUSY[31][0] , \ACCESS_BUSY[32][0] , 
        \ACCESS_BUSY[33][0] , \ACCESS_BUSY[34][0] , 
        \ACCESS_BUSY[35][0] , \ACCESS_BUSY[36][0] , 
        \ACCESS_BUSY[37][0] , \ACCESS_BUSY[38][0] , 
        \ACCESS_BUSY[39][0] , \ACCESS_BUSY[40][0] , 
        \ACCESS_BUSY[41][0] , \ACCESS_BUSY[42][0] , 
        \ACCESS_BUSY[43][0] , \ACCESS_BUSY[44][0] , 
        \ACCESS_BUSY[45][0] , \ACCESS_BUSY[46][0] , 
        \ACCESS_BUSY[47][0] , \ACCESS_BUSY[48][0] , 
        \ACCESS_BUSY[49][0] , \ACCESS_BUSY[50][0] , 
        \ACCESS_BUSY[51][0] , \ACCESS_BUSY[52][0] , 
        \ACCESS_BUSY[53][0] , \ACCESS_BUSY[54][0] , 
        \ACCESS_BUSY[55][0] , \ACCESS_BUSY[56][0] , 
        \ACCESS_BUSY[57][0] , \ACCESS_BUSY[58][0] , 
        \ACCESS_BUSY[59][0] , \ACCESS_BUSY[60][0] , 
        \ACCESS_BUSY[61][0] , \ACCESS_BUSY[62][0] , 
        \ACCESS_BUSY[63][0] , \ACCESS_BUSY[64][0] , 
        \ACCESS_BUSY[65][0] , \ACCESS_BUSY[66][0] , 
        \ACCESS_BUSY[67][0] , \ACCESS_BUSY[68][0] , 
        \ACCESS_BUSY[69][0] , \ACCESS_BUSY[70][0] , 
        \ACCESS_BUSY[71][0] , \ACCESS_BUSY[72][0] , 
        \ACCESS_BUSY[73][0] , \ACCESS_BUSY[74][0] , 
        \ACCESS_BUSY[75][0] , \ACCESS_BUSY[76][0] , 
        \ACCESS_BUSY[77][0] , \ACCESS_BUSY[78][0] , 
        \ACCESS_BUSY[79][0] , \ACCESS_BUSY[80][0] , 
        \ACCESS_BUSY[81][0] , \ACCESS_BUSY[82][0] , 
        \ACCESS_BUSY[83][0] , \ACCESS_BUSY[84][0] , 
        \ACCESS_BUSY[85][0] , \ACCESS_BUSY[86][0] , 
        \ACCESS_BUSY[87][0] , \ACCESS_BUSY[88][0] , 
        \ACCESS_BUSY[89][0] , \ACCESS_BUSY[90][0] , 
        \ACCESS_BUSY[91][0] , \ACCESS_BUSY[92][0] , 
        \ACCESS_BUSY[93][0] , \ACCESS_BUSY[94][0] , 
        \ACCESS_BUSY[95][0] , \ACCESS_BUSY[96][0] , 
        \ACCESS_BUSY[97][0] , \ACCESS_BUSY[98][0] , 
        \ACCESS_BUSY[99][0] , \ACCESS_BUSY[100][0] , 
        \ACCESS_BUSY[101][0] , \ACCESS_BUSY[102][0] , 
        \ACCESS_BUSY[103][0] , \ACCESS_BUSY[104][0] , 
        \ACCESS_BUSY[105][0] , \ACCESS_BUSY[106][0] , 
        \ACCESS_BUSY[107][0] , \ACCESS_BUSY[108][0] , 
        \ACCESS_BUSY[109][0] , \ACCESS_BUSY[110][0] , 
        \ACCESS_BUSY[111][0] , \ACCESS_BUSY[112][0] , 
        \ACCESS_BUSY[113][0] , \ACCESS_BUSY[114][0] , 
        \ACCESS_BUSY[115][0] , \ACCESS_BUSY[116][0] , 
        \ACCESS_BUSY[117][0] , \ACCESS_BUSY[118][0] , 
        \ACCESS_BUSY[119][0] , \ACCESS_BUSY[120][0] , 
        \ACCESS_BUSY[121][0] , \ACCESS_BUSY[122][0] , 
        \ACCESS_BUSY[123][0] , \ACCESS_BUSY[124][0] , 
        \ACCESS_BUSY[125][0] , \ACCESS_BUSY[126][0] , 
        \ACCESS_BUSY[127][0] , CFG3_16_Y, CFG3_15_Y, CFG3_0_Y, 
        CFG3_19_Y, CFG3_18_Y, CFG3_11_Y, CFG3_1_Y, CFG3_21_Y, CFG3_2_Y, 
        CFG3_20_Y, CFG3_9_Y, CFG3_3_Y, OR4_898_Y, OR4_809_Y, 
        OR4_1119_Y, OR4_1242_Y, OR4_1063_Y, OR4_506_Y, OR4_1071_Y, 
        OR4_455_Y, OR4_1089_Y, OR4_921_Y, OR4_1477_Y, OR4_292_Y, 
        OR4_1253_Y, OR4_1558_Y, OR4_999_Y, OR4_232_Y, OR4_1015_Y, 
        OR4_1284_Y, OR4_1487_Y, OR4_854_Y, OR4_1397_Y, OR4_209_Y, 
        OR4_1159_Y, OR4_1489_Y, OR4_918_Y, OR4_137_Y, OR4_943_Y, 
        OR4_1199_Y, OR4_1407_Y, OR4_1152_Y, OR4_70_Y, OR4_526_Y, 
        OR4_1495_Y, OR4_147_Y, OR4_1244_Y, OR4_469_Y, OR4_1258_Y, 
        OR4_1519_Y, OR4_74_Y, OR4_1275_Y, OR4_174_Y, OR2_17_Y, 
        OR4_215_Y, OR4_988_Y, OR4_1421_Y, OR4_1563_Y, OR4_358_Y, 
        OR4_1248_Y, OR4_247_Y, OR4_1012_Y, OR4_767_Y, OR4_1474_Y, 
        OR4_373_Y, OR4_1409_Y, OR4_4_Y, OR4_591_Y, OR4_1384_Y, 
        OR4_1635_Y, OR4_1129_Y, OR4_878_Y, OR4_596_Y, OR4_615_Y, 
        OR4_1143_Y, OR4_558_Y, OR4_791_Y, OR4_1380_Y, OR4_537_Y, 
        OR4_782_Y, OR4_300_Y, OR4_25_Y, OR4_1390_Y, OR4_1020_Y, 
        OR4_1572_Y, OR4_959_Y, OR4_1209_Y, OR4_142_Y, OR4_934_Y, 
        OR4_1192_Y, OR4_703_Y, OR4_447_Y, OR4_148_Y, OR4_1166_Y, 
        OR4_90_Y, OR2_26_Y, OR4_84_Y, OR4_454_Y, OR4_1185_Y, OR4_572_Y, 
        OR4_1587_Y, OR4_1235_Y, OR4_1603_Y, OR4_702_Y, OR4_689_Y, 
        OR4_508_Y, OR4_485_Y, OR4_152_Y, OR4_590_Y, OR4_416_Y, 
        OR4_1457_Y, OR4_344_Y, OR4_1478_Y, OR4_964_Y, OR4_1008_Y, 
        OR4_874_Y, OR4_853_Y, OR4_538_Y, OR4_952_Y, OR4_778_Y, 
        OR4_173_Y, OR4_696_Y, OR4_208_Y, OR4_1341_Y, OR4_1404_Y, 
        OR4_1617_Y, OR4_1596_Y, OR4_1270_Y, OR4_67_Y, OR4_1520_Y, 
        OR4_914_Y, OR4_1454_Y, OR4_936_Y, OR4_450_Y, OR4_504_Y, 
        OR4_981_Y, OR4_958_Y, OR2_18_Y, OR4_1383_Y, OR4_941_Y, 
        OR4_890_Y, OR4_827_Y, OR4_291_Y, OR4_1591_Y, OR4_1566_Y, 
        OR4_925_Y, OR4_653_Y, OR4_151_Y, OR4_126_Y, OR4_1469_Y, 
        OR4_249_Y, OR4_72_Y, OR4_1100_Y, OR4_1630_Y, OR4_1118_Y, 
        OR4_627_Y, OR4_677_Y, OR4_1376_Y, OR4_1349_Y, OR4_1014_Y, 
        OR4_1468_Y, OR4_1274_Y, OR4_668_Y, OR4_1190_Y, OR4_695_Y, 
        OR4_206_Y, OR4_257_Y, OR4_1318_Y, OR4_1283_Y, OR4_963_Y, 
        OR4_1406_Y, OR4_1214_Y, OR4_614_Y, OR4_1126_Y, OR4_636_Y, 
        OR4_128_Y, OR4_193_Y, OR4_1254_Y, OR4_1228_Y, OR2_25_Y, 
        OR4_398_Y, OR4_847_Y, OR4_718_Y, OR4_843_Y, OR4_496_Y, 
        OR4_1018_Y, OR4_1450_Y, OR4_553_Y, OR4_665_Y, OR4_430_Y, 
        OR4_957_Y, OR4_1423_Y, OR4_748_Y, OR4_1051_Y, OR4_513_Y, 
        OR4_1367_Y, OR4_535_Y, OR4_781_Y, OR4_967_Y, OR4_884_Y, 
        OR4_1424_Y, OR4_238_Y, OR4_1197_Y, OR4_1510_Y, OR4_955_Y, 
        OR4_179_Y, OR4_974_Y, OR4_1234_Y, OR4_1436_Y, OR4_754_Y, 
        OR4_1293_Y, OR4_108_Y, OR4_1070_Y, OR4_1396_Y, OR4_830_Y, 
        OR4_60_Y, OR4_856_Y, OR4_1108_Y, OR4_1305_Y, OR4_879_Y, 
        OR4_1422_Y, OR2_6_Y, OR4_314_Y, OR4_85_Y, OR4_962_Y, 
        OR4_1187_Y, OR4_1444_Y, OR4_1088_Y, OR4_821_Y, OR4_904_Y, 
        OR4_855_Y, OR4_717_Y, OR4_693_Y, OR4_380_Y, OR4_799_Y, 
        OR4_626_Y, OR4_19_Y, OR4_554_Y, OR4_49_Y, OR4_1178_Y, 
        OR4_1238_Y, OR4_511_Y, OR4_488_Y, OR4_154_Y, OR4_594_Y, 
        OR4_417_Y, OR4_1458_Y, OR4_346_Y, OR4_1480_Y, OR4_965_Y, 
        OR4_1010_Y, OR4_1400_Y, OR4_1374_Y, OR4_1037_Y, OR4_1486_Y, 
        OR4_1301_Y, OR4_688_Y, OR4_1213_Y, OR4_716_Y, OR4_222_Y, 
        OR4_276_Y, OR4_1618_Y, OR4_1600_Y, OR2_31_Y, OR4_818_Y, 
        OR4_1002_Y, OR4_608_Y, OR4_1219_Y, OR4_252_Y, OR4_356_Y, 
        OR4_877_Y, OR4_343_Y, OR4_1075_Y, OR4_858_Y, OR4_1403_Y, 
        OR4_212_Y, OR4_1162_Y, OR4_1492_Y, OR4_928_Y, OR4_141_Y, 
        OR4_948_Y, OR4_1206_Y, OR4_1410_Y, OR4_1035_Y, OR4_1585_Y, 
        OR4_407_Y, OR4_1377_Y, OR4_40_Y, OR4_1117_Y, OR4_361_Y, 
        OR4_1135_Y, OR4_1414_Y, OR4_1595_Y, OR4_643_Y, OR4_1168_Y, 
        OR4_1633_Y, OR4_961_Y, OR4_1271_Y, OR4_723_Y, OR4_1577_Y, 
        OR4_740_Y, OR4_990_Y, OR4_1177_Y, OR4_1255_Y, OR4_146_Y, 
        OR2_15_Y, OR4_625_Y, OR4_1514_Y, OR4_163_Y, OR4_261_Y, 
        OR4_1425_Y, OR4_922_Y, OR4_1006_Y, OR4_1315_Y, OR4_265_Y, 
        OR4_248_Y, OR4_783_Y, OR4_177_Y, OR4_429_Y, OR4_996_Y, 
        OR4_145_Y, OR4_420_Y, OR4_1552_Y, OR4_1296_Y, OR4_1000_Y, 
        OR4_1121_Y, OR4_37_Y, OR4_1057_Y, OR4_1322_Y, OR4_263_Y, 
        OR4_1031_Y, OR4_1306_Y, OR4_802_Y, OR4_552_Y, OR4_266_Y, 
        OR4_1432_Y, OR4_341_Y, OR4_1360_Y, OR4_1607_Y, OR4_551_Y, 
        OR4_1337_Y, OR4_1597_Y, OR4_1091_Y, OR4_834_Y, OR4_559_Y, 
        OR4_1504_Y, OR4_418_Y, OR2_35_Y, OR4_390_Y, OR4_20_Y, 
        OR4_1543_Y, OR4_1266_Y, OR4_1030_Y, OR4_1588_Y, OR4_656_Y, 
        OR4_1329_Y, OR4_733_Y, OR4_1637_Y, OR4_546_Y, OR4_1571_Y, 
        OR4_180_Y, OR4_759_Y, OR4_1542_Y, OR4_166_Y, OR4_1321_Y, 
        OR4_1042_Y, OR4_764_Y, OR4_1277_Y, OR4_184_Y, OR4_1212_Y, 
        OR4_1473_Y, OR4_408_Y, OR4_1186_Y, OR4_1465_Y, OR4_951_Y, 
        OR4_687_Y, OR4_411_Y, OR4_1157_Y, OR4_73_Y, OR4_1093_Y, 
        OR4_1351_Y, OR4_298_Y, OR4_1072_Y, OR4_1338_Y, OR4_844_Y, 
        OR4_585_Y, OR4_303_Y, OR4_889_Y, OR4_1437_Y, OR2_23_Y, 
        OR4_269_Y, OR4_1553_Y, OR4_1029_Y, OR4_1358_Y, OR4_741_Y, 
        OR4_1297_Y, OR4_1155_Y, OR4_499_Y, OR4_267_Y, OR4_321_Y, 
        OR4_836_Y, OR4_1289_Y, OR4_622_Y, OR4_923_Y, OR4_382_Y, 
        OR4_1230_Y, OR4_404_Y, OR4_657_Y, OR4_846_Y, OR4_1599_Y, 
        OR4_500_Y, OR4_942_Y, OR4_288_Y, OR4_592_Y, OR4_36_Y, 
        OR4_895_Y, OR4_59_Y, OR4_327_Y, OR4_510_Y, OR4_1076_Y, 
        OR4_1619_Y, OR4_437_Y, OR4_1411_Y, OR4_76_Y, OR4_1145_Y, 
        OR4_379_Y, OR4_1163_Y, OR4_1443_Y, OR4_1628_Y, OR4_1401_Y, 
        OR4_296_Y, OR2_21_Y, OR4_389_Y, OR4_319_Y, OR4_342_Y, 
        OR4_1470_Y, OR4_929_Y, OR4_1208_Y, OR4_1203_Y, OR4_1488_Y, 
        OR4_779_Y, OR4_798_Y, OR4_780_Y, OR4_468_Y, OR4_892_Y, 
        OR4_710_Y, OR4_112_Y, OR4_630_Y, OR4_124_Y, OR4_1269_Y, 
        OR4_1330_Y, OR4_721_Y, OR4_699_Y, OR4_385_Y, OR4_801_Y, 
        OR4_629_Y, OR4_22_Y, OR4_557_Y, OR4_54_Y, OR4_1181_Y, 
        OR4_1241_Y, OR4_747_Y, OR4_728_Y, OR4_414_Y, OR4_831_Y, 
        OR4_659_Y, OR4_61_Y, OR4_582_Y, OR4_83_Y, OR4_1215_Y, 
        OR4_1267_Y, OR4_243_Y, OR4_220_Y, OR2_39_Y, OR4_1038_Y, 
        OR4_991_Y, OR4_772_Y, OR4_38_Y, OR4_1347_Y, OR4_670_Y, 
        OR4_1005_Y, OR4_196_Y, OR4_322_Y, OR4_663_Y, OR4_1200_Y, 
        OR4_603_Y, OR4_849_Y, OR4_1433_Y, OR4_583_Y, OR4_832_Y, 
        OR4_355_Y, OR4_82_Y, OR4_1440_Y, OR4_617_Y, OR4_1147_Y, 
        OR4_560_Y, OR4_793_Y, OR4_1386_Y, OR4_539_Y, OR4_785_Y, 
        OR4_304_Y, OR4_29_Y, OR4_1392_Y, OR4_393_Y, OR4_919_Y, 
        OR4_336_Y, OR4_574_Y, OR4_1136_Y, OR4_317_Y, OR4_565_Y, 
        OR4_68_Y, OR4_1447_Y, OR4_1137_Y, OR4_1290_Y, OR4_198_Y, 
        OR2_29_Y, OR4_360_Y, OR4_1124_Y, OR4_1544_Y, OR4_66_Y, 
        OR4_486_Y, OR4_1393_Y, OR4_386_Y, OR4_1148_Y, OR4_905_Y, 
        OR4_931_Y, OR4_909_Y, OR4_62_Y, OR4_528_Y, OR4_826_Y, 
        OR4_1065_Y, OR4_883_Y, OR4_522_Y, OR4_363_Y, OR4_481_Y, 
        OR4_94_Y, OR4_65_Y, OR4_845_Y, OR4_1316_Y, OR4_1621_Y, 
        OR4_228_Y, OR4_30_Y, OR4_1308_Y, OR4_1127_Y, OR4_1260_Y, 
        OR4_512_Y, OR4_480_Y, OR4_1256_Y, OR4_92_Y, OR4_406_Y, 
        OR4_641_Y, OR4_452_Y, OR4_88_Y, OR4_1546_Y, OR4_43_Y, 
        OR4_654_Y, OR4_623_Y, OR2_34_Y, OR4_1288_Y, OR4_440_Y, 
        OR4_1059_Y, OR4_605_Y, OR4_311_Y, OR4_1243_Y, OR4_1323_Y, 
        OR4_516_Y, OR4_1441_Y, OR4_906_Y, OR4_1461_Y, OR4_841_Y, 
        OR4_1084_Y, OR4_26_Y, OR4_815_Y, OR4_1067_Y, OR4_586_Y, 
        OR4_333_Y, OR4_31_Y, OR4_50_Y, OR4_598_Y, OR4_1623_Y, 
        OR4_235_Y, OR4_804_Y, OR4_1604_Y, OR4_224_Y, OR4_1370_Y, 
        OR4_1094_Y, OR4_810_Y, OR4_681_Y, OR4_1224_Y, OR4_619_Y, 
        OR4_869_Y, OR4_1459_Y, OR4_601_Y, OR4_859_Y, OR4_370_Y, 
        OR4_104_Y, OR4_1462_Y, OR4_226_Y, OR4_762_Y, OR2_2_Y, 
        OR4_953_Y, OR4_1499_Y, OR4_1032_Y, OR4_800_Y, OR4_1569_Y, 
        OR4_242_Y, OR4_1193_Y, OR4_1004_Y, OR4_448_Y, OR4_986_Y, 
        OR4_1527_Y, OR4_362_Y, OR4_1326_Y, OR4_1627_Y, OR4_1061_Y, 
        OR4_302_Y, OR4_1086_Y, OR4_1352_Y, OR4_1533_Y, OR4_1526_Y, 
        OR4_431_Y, OR4_885_Y, OR4_217_Y, OR4_532_Y, OR4_1608_Y, 
        OR4_824_Y, OR4_1631_Y, OR4_254_Y, OR4_444_Y, OR4_1079_Y, 
        OR4_1620_Y, OR4_439_Y, OR4_1413_Y, OR4_79_Y, OR4_1146_Y, 
        OR4_381_Y, OR4_1164_Y, OR4_1446_Y, OR4_1629_Y, OR4_842_Y, 
        OR4_1389_Y, OR2_4_Y, OR4_766_Y, OR4_10_Y, OR4_323_Y, OR4_395_Y, 
        OR4_1549_Y, OR4_1058_Y, OR4_1139_Y, OR4_1456_Y, OR4_403_Y, 
        OR4_1359_Y, OR4_1332_Y, OR4_476_Y, OR4_930_Y, OR4_1249_Y, 
        OR4_1496_Y, OR4_1302_Y, OR4_926_Y, OR4_770_Y, OR4_896_Y, 
        OR4_607_Y, OR4_581_Y, OR4_1363_Y, OR4_185_Y, OR4_507_Y, 
        OR4_742_Y, OR4_555_Y, OR4_183_Y, OR4_12_Y, OR4_132_Y, 
        OR4_900_Y, OR4_871_Y, OR4_9_Y, OR4_482_Y, OR4_788_Y, 
        OR4_1021_Y, OR4_839_Y, OR4_475_Y, OR4_325_Y, OR4_442_Y, 
        OR4_976_Y, OR4_947_Y, OR2_0_Y, OR4_527_Y, OR4_157_Y, OR4_47_Y, 
        OR4_1415_Y, OR4_1167_Y, OR4_91_Y, OR4_787_Y, OR4_1471_Y, 
        OR4_875_Y, OR4_1106_Y, OR4_1081_Y, OR4_230_Y, OR4_685_Y, 
        OR4_997_Y, OR4_1247_Y, OR4_1046_Y, OR4_683_Y, OR4_530_Y, 
        OR4_649_Y, OR4_751_Y, OR4_726_Y, OR4_1506_Y, OR4_352_Y, 
        OR4_648_Y, OR4_893_Y, OR4_692_Y, OR4_349_Y, OR4_161_Y, 
        OR4_301_Y, OR4_640_Y, OR4_610_Y, OR4_1408_Y, OR4_227_Y, 
        OR4_541_Y, OR4_776_Y, OR4_588_Y, OR4_218_Y, OR4_52_Y, 
        OR4_175_Y, OR4_369_Y, OR4_347_Y, OR2_27_Y, CFG3_13_Y, CFG3_8_Y, 
        CFG3_14_Y, CFG3_5_Y, CFG3_6_Y, CFG3_22_Y, CFG3_10_Y, CFG3_23_Y, 
        CFG3_12_Y, CFG3_4_Y, CFG3_17_Y, CFG3_7_Y, OR4_1331_Y, 
        OR4_1529_Y, OR4_1077_Y, OR4_866_Y, OR4_1502_Y, OR4_23_Y, 
        OR4_143_Y, OR4_33_Y, OR4_971_Y, OR4_1365_Y, OR4_268_Y, 
        OR4_711_Y, OR4_45_Y, OR4_368_Y, OR4_1451_Y, OR4_660_Y, 
        OR4_1472_Y, OR4_86_Y, OR4_274_Y, OR4_1567_Y, OR4_472_Y, 
        OR4_915_Y, OR4_259_Y, OR4_567_Y, OR4_5_Y, OR4_868_Y, OR4_24_Y, 
        OR4_293_Y, OR4_478_Y, OR4_1110_Y, OR4_11_Y, OR4_473_Y, 
        OR4_1449_Y, OR4_109_Y, OR4_1188_Y, OR4_422_Y, OR4_1210_Y, 
        OR4_1485_Y, OR4_17_Y, OR4_903_Y, OR4_1445_Y, OR2_8_Y, 
        OR4_1171_Y, OR4_1128_Y, OR4_907_Y, OR4_170_Y, OR4_1491_Y, 
        OR4_806_Y, OR4_1138_Y, OR4_345_Y, OR4_446_Y, OR4_127_Y, 
        OR4_110_Y, OR4_897_Y, OR4_1361_Y, OR4_32_Y, OR4_281_Y, 
        OR4_89_Y, OR4_1355_Y, OR4_1173_Y, OR4_1324_Y, OR4_98_Y, 
        OR4_69_Y, OR4_850_Y, OR4_1319_Y, OR4_1626_Y, OR4_231_Y, 
        OR4_34_Y, OR4_1314_Y, OR4_1130_Y, OR4_1264_Y, OR4_1501_Y, 
        OR4_1479_Y, OR4_616_Y, OR4_1073_Y, OR4_1405_Y, OR4_1636_Y, 
        OR4_1453_Y, OR4_1066_Y, OR4_910_Y, OR4_1023_Y, OR4_768_Y, 
        OR4_732_Y, OR2_37_Y, OR4_1435_Y, OR4_576_Y, OR4_1196_Y, 
        OR4_738_Y, OR4_436_Y, OR4_1387_Y, OR4_1463_Y, OR4_646_Y, 
        OR4_1568_Y, OR4_383_Y, OR4_364_Y, OR4_1125_Y, OR4_1602_Y, 
        OR4_278_Y, OR4_524_Y, OR4_337_Y, OR4_1598_Y, OR4_1438_Y, 
        OR4_1548_Y, OR4_1149_Y, OR4_1122_Y, OR4_286_Y, OR4_743_Y, 
        OR4_1048_Y, OR4_1298_Y, OR4_1102_Y, OR4_734_Y, OR4_578_Y, 
        OR4_697_Y, OR4_149_Y, OR4_122_Y, OR4_912_Y, OR4_1385_Y, 
        OR4_56_Y, OR4_307_Y, OR4_105_Y, OR4_1379_Y, OR4_1201_Y, 
        OR4_1336_Y, OR4_1335_Y, OR4_1309_Y, OR2_10_Y, OR4_1428_Y, 
        OR4_851_Y, OR4_8_Y, OR4_722_Y, OR4_1142_Y, OR4_1503_Y, 
        OR4_42_Y, OR4_1236_Y, OR4_1282_Y, OR4_1025_Y, OR4_1576_Y, 
        OR4_969_Y, OR4_1216_Y, OR4_153_Y, OR4_945_Y, OR4_1202_Y, 
        OR4_709_Y, OR4_459_Y, OR4_159_Y, OR4_470_Y, OR4_998_Y, 
        OR4_405_Y, OR4_644_Y, OR4_1222_Y, OR4_377_Y, OR4_632_Y, 
        OR4_129_Y, OR4_1515_Y, OR4_1225_Y, OR4_1261_Y, OR4_164_Y, 
        OR4_1191_Y, OR4_1460_Y, OR4_392_Y, OR4_1161_Y, OR4_1442_Y, 
        OR4_933_Y, OR4_672_Y, OR4_399_Y, OR4_353_Y, OR4_882_Y, OR2_9_Y, 
        OR4_219_Y, OR4_529_Y, OR4_939_Y, OR4_1259_Y, OR4_521_Y, 
        OR4_1448_Y, OR4_908_Y, OR4_365_Y, OR4_852_Y, OR4_264_Y, 
        OR4_789_Y, OR4_1246_Y, OR4_584_Y, OR4_887_Y, OR4_350_Y, 
        OR4_1182_Y, OR4_366_Y, OR4_611_Y, OR4_792_Y, OR4_564_Y, 
        OR4_1087_Y, OR4_1541_Y, OR4_881_Y, OR4_1174_Y, OR4_633_Y, 
        OR4_1497_Y, OR4_655_Y, OR4_911_Y, OR4_1092_Y, OR4_977_Y, 
        OR4_1518_Y, OR4_351_Y, OR4_1311_Y, OR4_1614_Y, OR4_1054_Y, 
        OR4_289_Y, OR4_1074_Y, OR4_1339_Y, OR4_1522_Y, OR4_1303_Y, 
        OR4_204_Y, OR2_19_Y, OR4_724_Y, OR4_1509_Y, OR4_297_Y, 
        OR4_445_Y, OR4_860_Y, OR4_117_Y, OR4_758_Y, OR4_1532_Y, 
        OR4_1272_Y, OR4_1132_Y, OR4_1112_Y, OR4_796_Y, OR4_1226_Y, 
        OR4_1044_Y, OR4_453_Y, OR4_968_Y, OR4_477_Y, OR4_1615_Y, 
        OR4_21_Y, OR4_305_Y, OR4_277_Y, OR4_1593_Y, OR4_384_Y, 
        OR4_211_Y, OR4_1231_Y, OR4_118_Y, OR4_1257_Y, OR4_763_Y, 
        OR4_812_Y, OR4_708_Y, OR4_684_Y, OR4_374_Y, OR4_790_Y, 
        OR4_620_Y, OR4_13_Y, OR4_545_Y, OR4_41_Y, OR4_1165_Y, 
        OR4_1227_Y, OR4_862_Y, OR4_837_Y, OR2_12_Y, OR4_1354_Y, 
        OR4_1539_Y, OR4_1016_Y, OR4_1340_Y, OR4_1292_Y, OR4_1280_Y, 
        OR4_1169_Y, OR4_1582_Y, OR4_251_Y, OR4_1399_Y, OR4_294_Y, 
        OR4_739_Y, OR4_78_Y, OR4_387_Y, OR4_1476_Y, OR4_682_Y, 
        OR4_1494_Y, OR4_107_Y, OR4_309_Y, OR4_1578_Y, OR4_487_Y, 
        OR4_927_Y, OR4_271_Y, OR4_580_Y, OR4_15_Y, OR4_880_Y, OR4_39_Y, 
        OR4_318_Y, OR4_495_Y, OR4_1056_Y, OR4_1606_Y, OR4_425_Y, 
        OR4_1398_Y, OR4_64_Y, OR4_1133_Y, OR4_371_Y, OR4_1151_Y, 
        OR4_1430_Y, OR4_1611_Y, OR4_1382_Y, OR4_282_Y, OR2_20_Y, 
        OR4_1195_Y, OR4_1574_Y, OR4_675_Y, OR4_55_Y, OR4_1064_Y, 
        OR4_727_Y, OR4_1085_Y, OR4_197_Y, OR4_182_Y, OR4_820_Y, 
        OR4_1366_Y, OR4_753_Y, OR4_993_Y, OR4_1581_Y, OR4_729_Y, 
        OR4_984_Y, OR4_503_Y, OR4_237_Y, OR4_1586_Y, OR4_1184_Y, 
        OR4_102_Y, OR4_1115_Y, OR4_1378_Y, OR4_328_Y, OR4_1101_Y, 
        OR4_1364_Y, OR4_870_Y, OR4_606_Y, OR4_331_Y, OR4_313_Y, 
        OR4_838_Y, OR4_234_Y, OR4_484_Y, OR4_1050_Y, OR4_214_Y, 
        OR4_471_Y, OR4_1610_Y, OR4_1350_Y, OR4_1055_Y, OR4_1313_Y, 
        OR4_216_Y, OR2_30_Y, OR4_865_Y, OR4_441_Y, OR4_375_Y, 
        OR4_335_Y, OR4_1416_Y, OR4_1069_Y, OR4_1045_Y, OR4_426_Y, 
        OR4_130_Y, OR4_489_Y, OR4_1009_Y, OR4_421_Y, OR4_661_Y, 
        OR4_1239_Y, OR4_401_Y, OR4_651_Y, OR4_144_Y, OR4_1528_Y, 
        OR4_1245_Y, OR4_51_Y, OR4_599_Y, OR4_1624_Y, OR4_236_Y, 
        OR4_805_Y, OR4_1605_Y, OR4_225_Y, OR4_1371_Y, OR4_1095_Y, 
        OR4_811_Y, OR4_1632_Y, OR4_540_Y, OR4_1564_Y, OR4_169_Y, 
        OR4_750_Y, OR4_1536_Y, OR4_155_Y, OR4_1310_Y, OR4_1027_Y, 
        OR4_752_Y, OR4_1573_Y, OR4_483_Y, OR2_36_Y, OR4_1131_Y, 
        OR4_397_Y, OR4_676_Y, OR4_769_Y, OR4_306_Y, OR4_1455_Y, 
        OR4_1524_Y, OR4_181_Y, OR4_773_Y, OR4_1561_Y, OR4_1535_Y, 
        OR4_1217_Y, OR4_7_Y, OR4_1484_Y, OR4_872_Y, OR4_1402_Y, 
        OR4_894_Y, OR4_402_Y, OR4_449_Y, OR4_807_Y, OR4_786_Y, 
        OR4_474_Y, OR4_902_Y, OR4_720_Y, OR4_114_Y, OR4_638_Y, 
        OR4_131_Y, OR4_1276_Y, OR4_1333_Y, OR4_1097_Y, OR4_1080_Y, 
        OR4_761_Y, OR4_1179_Y, OR4_1003_Y, OR4_413_Y, OR4_920_Y, 
        OR4_438_Y, OR4_1570_Y, OR4_1625_Y, OR4_1175_Y, OR4_1153_Y, 
        OR2_24_Y, OR4_1551_Y, OR4_979_Y, OR4_135_Y, OR4_861_Y, 
        OR4_1291_Y, OR4_1638_Y, OR4_176_Y, OR4_1381_Y, OR4_1429_Y, 
        OR4_517_Y, OR4_490_Y, OR4_1263_Y, OR4_97_Y, OR4_409_Y, 
        OR4_647_Y, OR4_461_Y, OR4_93_Y, OR4_1555_Y, OR4_48_Y, 
        OR4_1575_Y, OR4_1540_Y, OR4_686_Y, OR4_1144_Y, OR4_1481_Y, 
        OR4_80_Y, OR4_1517_Y, OR4_1140_Y, OR4_982_Y, OR4_1109_Y, 
        OR4_735_Y, OR4_704_Y, OR4_1498_Y, OR4_334_Y, OR4_631_Y, 
        OR4_876_Y, OR4_678_Y, OR4_329_Y, OR4_138_Y, OR4_283_Y, 
        OR4_1464_Y, OR4_1426_Y, OR2_14_Y, OR4_899_Y, OR4_544_Y, 
        OR4_428_Y, OR4_133_Y, OR4_1550_Y, OR4_467_Y, OR4_1156_Y, 
        OR4_202_Y, OR4_1250_Y, OR4_1327_Y, OR4_1295_Y, OR4_972_Y, 
        OR4_1412_Y, OR4_1223_Y, OR4_621_Y, OR4_1134_Y, OR4_645_Y, 
        OR4_136_Y, OR4_207_Y, OR4_954_Y, OR4_932_Y, OR4_618_Y, 
        OR4_1034_Y, OR4_873_Y, OR4_272_Y, OR4_784_Y, OR4_299_Y, 
        OR4_1439_Y, OR4_1490_Y, OR4_848_Y, OR4_823_Y, OR4_514_Y, 
        OR4_924_Y, OR4_755_Y, OR4_139_Y, OR4_669_Y, OR4_172_Y, 
        OR4_1325_Y, OR4_1373_Y, OR4_573_Y, OR4_549_Y, OR2_5_Y, 
        OR4_1431_Y, OR4_1198_Y, OR4_462_Y, OR4_679_Y, OR4_917_Y, 
        OR4_587_Y, OR4_326_Y, OR4_394_Y, OR4_354_Y, OR4_1026_Y, 
        OR4_1580_Y, OR4_970_Y, OR4_1218_Y, OR4_156_Y, OR4_946_Y, 
        OR4_1204_Y, OR4_712_Y, OR4_460_Y, OR4_162_Y, OR4_822_Y, 
        OR4_1369_Y, OR4_756_Y, OR4_994_Y, OR4_1583_Y, OR4_730_Y, 
        OR4_985_Y, OR4_505_Y, OR4_239_Y, OR4_1589_Y, OR4_75_Y, 
        OR4_613_Y, OR4_1_Y, OR4_260_Y, OR4_825_Y, OR4_1622_Y, 
        OR4_244_Y, OR4_1394_Y, OR4_1113_Y, OR4_833_Y, OR4_316_Y, 
        OR4_840_Y, OR2_7_Y, OR4_1557_Y, OR4_1512_Y, OR4_1279_Y, 
        OR4_556_Y, OR4_223_Y, OR4_1176_Y, OR4_1523_Y, OR4_701_Y, 
        OR4_814_Y, OR4_359_Y, OR4_339_Y, OR4_1639_Y, OR4_432_Y, 
        OR4_262_Y, OR4_1285_Y, OR4_168_Y, OR4_1320_Y, OR4_808_Y, 
        OR4_867_Y, OR4_315_Y, OR4_285_Y, OR4_1601_Y, OR4_391_Y, 
        OR4_213_Y, OR4_1240_Y, OR4_121_Y, OR4_1262_Y, OR4_771_Y, 
        OR4_819_Y, OR4_71_Y, OR4_44_Y, OR4_1368_Y, OR4_140_Y, 
        OR4_1616_Y, OR4_1001_Y, OR4_1530_Y, OR4_1022_Y, OR4_542_Y, 
        OR4_595_Y, OR4_966_Y, OR4_944_Y, OR2_16_Y, OR4_388_Y, 
        OR4_1154_Y, OR4_63_Y, OR4_295_Y, OR4_229_Y, OR4_757_Y, 
        OR4_400_Y, OR4_396_Y, OR4_338_Y, OR4_424_Y, OR4_950_Y, 
        OR4_1417_Y, OR4_737_Y, OR4_1036_Y, OR4_502_Y, OR4_1357_Y, 
        OR4_523_Y, OR4_775_Y, OR4_956_Y, OR4_1194_Y, OR4_106_Y, 
        OR4_562_Y, OR4_1521_Y, OR4_199_Y, OR4_1278_Y, OR4_509_Y, 
        OR4_1304_Y, OR4_1556_Y, OR4_111_Y, OR4_100_Y, OR4_628_Y, 
        OR4_1082_Y, OR4_423_Y, OR4_725_Y, OR4_167_Y, OR4_1017_Y, 
        OR4_191_Y, OR4_456_Y, OR4_635_Y, OR4_340_Y, OR4_863_Y, 
        OR2_33_Y, OR4_158_Y, OR4_940_Y, OR4_1579_Y, OR4_1111_Y, 
        OR4_803_Y, OR4_115_Y, OR4_188_Y, OR4_1011_Y, OR4_324_Y, 
        OR4_589_Y, OR4_571_Y, OR4_246_Y, OR4_666_Y, OR4_501_Y, 
        OR4_1525_Y, OR4_419_Y, OR4_1547_Y, OR4_1047_Y, OR4_1105_Y, 
        OR4_1375_Y, OR4_1348_Y, OR4_1013_Y, OR4_1467_Y, OR4_1273_Y, 
        OR4_667_Y, OR4_1189_Y, OR4_694_Y, OR4_205_Y, OR4_256_Y, 
        OR4_372_Y, OR4_357_Y, OR4_18_Y, OR4_458_Y, OR4_279_Y, 
        OR4_1317_Y, OR4_195_Y, OR4_1334_Y, OR4_829_Y, OR4_888_Y, 
        OR4_1534_Y, OR4_1516_Y, OR2_28_Y, OR4_1505_Y, OR4_1434_Y, 
        OR4_1466_Y, OR4_937_Y, OR4_427_Y, OR4_700_Y, OR4_691_Y, 
        OR4_960_Y, OR4_275_Y, OR4_1114_Y, OR4_27_Y, OR4_1052_Y, 
        OR4_1312_Y, OR4_253_Y, OR4_1024_Y, OR4_1294_Y, OR4_794_Y, 
        OR4_543_Y, OR4_258_Y, OR4_1028_Y, OR4_1584_Y, OR4_973_Y, 
        OR4_1220_Y, OR4_160_Y, OR4_949_Y, OR4_1207_Y, OR4_714_Y, 
        OR4_463_Y, OR4_165_Y, OR4_1060_Y, OR4_1612_Y, OR4_995_Y, 
        OR4_1251_Y, OR4_194_Y, OR4_975_Y, OR4_1237_Y, OR4_745_Y, 
        OR4_491_Y, OR4_201_Y, OR4_570_Y, OR4_1098_Y, OR2_11_Y, 
        OR4_1342_Y, OR4_77_Y, OR4_813_Y, OR4_186_Y, OR4_1205_Y, 
        OR4_864_Y, OR4_1221_Y, OR4_348_Y, OR4_332_Y, OR4_308_Y, 
        OR4_270_Y, OR4_1041_Y, OR4_1511_Y, OR4_189_Y, OR4_433_Y, 
        OR4_240_Y, OR4_1507_Y, OR4_1344_Y, OR4_1482_Y, OR4_664_Y, 
        OR4_634_Y, OR4_1427_Y, OR4_250_Y, OR4_566_Y, OR4_795_Y, 
        OR4_609_Y, OR4_245_Y, OR4_81_Y, OR4_210_Y, OR4_1418_Y, 
        OR4_1388_Y, OR4_536_Y, OR4_983_Y, OR4_1307_Y, OR4_1538_Y, 
        OR4_1353_Y, OR4_980_Y, OR4_817_Y, OR4_938_Y, OR4_777_Y, 
        OR4_749_Y, OR2_38_Y, OR4_1252_Y, OR4_330_Y, OR4_534_Y, 
        OR4_707_Y, OR4_192_Y, OR4_497_Y, OR4_203_Y, OR4_1040_Y, 
        OR4_123_Y, OR4_1287_Y, OR4_187_Y, OR4_642_Y, OR4_1613_Y, 
        OR4_290_Y, OR4_1372_Y, OR4_593_Y, OR4_1395_Y, OR4_3_Y, 
        OR4_200_Y, OR4_367_Y, OR4_891_Y, OR4_1345_Y, OR4_671_Y, 
        OR4_978_Y, OR4_434_Y, OR4_1286_Y, OR4_457_Y, OR4_706_Y, 
        OR4_901_Y, OR4_569_Y, OR4_1090_Y, OR4_1545_Y, OR4_886_Y, 
        OR4_1183_Y, OR4_637_Y, OR4_1500_Y, OR4_658_Y, OR4_913_Y, 
        OR4_1104_Y, OR4_746_Y, OR4_1281_Y, OR2_1_Y, OR4_989_Y, 
        OR4_577_Y, OR4_515_Y, OR4_465_Y, OR4_1537_Y, OR4_1211_Y, 
        OR4_1180_Y, OR4_563_Y, OR4_284_Y, OR4_1594_Y, OR4_1562_Y, 
        OR4_705_Y, OR4_1160_Y, OR4_1493_Y, OR4_96_Y, OR4_1531_Y, 
        OR4_1158_Y, OR4_992_Y, OR4_1120_Y, OR4_1150_Y, OR4_1123_Y, 
        OR4_287_Y, OR4_744_Y, OR4_1049_Y, OR4_1299_Y, OR4_1103_Y, 
        OR4_736_Y, OR4_579_Y, OR4_698_Y, OR4_1099_Y, OR4_1062_Y, 
        OR4_221_Y, OR4_680_Y, OR4_987_Y, OR4_1233_Y, OR4_1033_Y, 
        OR4_673_Y, OR4_518_Y, OR4_639_Y, OR4_1039_Y, OR4_1007_Y, 
        OR2_3_Y, OR4_1554_Y, OR4_1343_Y, OR4_597_Y, OR4_816_Y, 
        OR4_1053_Y, OR4_715_Y, OR4_451_Y, OR4_533_Y, OR4_479_Y, 
        OR4_519_Y, OR4_492_Y, OR4_1265_Y, OR4_101_Y, OR4_412_Y, 
        OR4_650_Y, OR4_464_Y, OR4_95_Y, OR4_1559_Y, OR4_53_Y, 
        OR4_312_Y, OR4_273_Y, OR4_1043_Y, OR4_1513_Y, OR4_190_Y, 
        OR4_435_Y, OR4_241_Y, OR4_1508_Y, OR4_1346_Y, OR4_1483_Y, 
        OR4_1170_Y, OR4_1141_Y, OR4_320_Y, OR4_765_Y, OR4_1068_Y, 
        OR4_1328_Y, OR4_1116_Y, OR4_760_Y, OR4_600_Y, OR4_719_Y, 
        OR4_1419_Y, OR4_1391_Y, OR2_13_Y, OR4_2_Y, OR4_1560_Y, 
        OR4_1590_Y, OR4_1078_Y, OR4_568_Y, OR4_835_Y, OR4_828_Y, 
        OR4_1096_Y, OR4_410_Y, OR4_602_Y, OR4_575_Y, OR4_1356_Y, 
        OR4_178_Y, OR4_498_Y, OR4_731_Y, OR4_547_Y, OR4_171_Y, OR4_6_Y, 
        OR4_125_Y, OR4_525_Y, OR4_494_Y, OR4_1268_Y, OR4_103_Y, 
        OR4_415_Y, OR4_652_Y, OR4_466_Y, OR4_99_Y, OR4_1565_Y, 
        OR4_57_Y, OR4_548_Y, OR4_520_Y, OR4_1300_Y, OR4_120_Y, 
        OR4_443_Y, OR4_674_Y, OR4_493_Y, OR4_116_Y, OR4_1592_Y, 
        OR4_87_Y, OR4_35_Y, OR4_0_Y, OR2_22_Y, OR4_310_Y, OR4_1362_Y, 
        OR4_531_Y, OR4_1229_Y, OR4_28_Y, OR4_378_Y, OR4_561_Y, 
        OR4_113_Y, OR4_150_Y, OR4_713_Y, OR4_690_Y, OR4_376_Y, 
        OR4_797_Y, OR4_624_Y, OR4_16_Y, OR4_550_Y, OR4_46_Y, 
        OR4_1172_Y, OR4_1232_Y, OR4_134_Y, OR4_119_Y, OR4_1452_Y, 
        OR4_233_Y, OR4_58_Y, OR4_1083_Y, OR4_1609_Y, OR4_1107_Y, 
        OR4_612_Y, OR4_662_Y, OR4_935_Y, OR4_916_Y, OR4_604_Y, 
        OR4_1019_Y, OR4_857_Y, OR4_255_Y, OR4_774_Y, OR4_280_Y, 
        OR4_1420_Y, OR4_1475_Y, OR4_14_Y, OR4_1634_Y, OR2_32_Y, VCC, 
        GND, ADLIB_VCC;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign ADLIB_VCC = VCC_power_net1;
    
    OR4 OR4_700 (.A(OR4_949_Y), .B(OR4_1207_Y), .C(OR4_714_Y), .D(
        OR4_463_Y), .Y(OR4_700_Y));
    OR4 OR4_399 (.A(\R_DATA_TEMPR72[24] ), .B(\R_DATA_TEMPR73[24] ), 
        .C(\R_DATA_TEMPR74[24] ), .D(\R_DATA_TEMPR75[24] ), .Y(
        OR4_399_Y));
    OR4 OR4_1188 (.A(\R_DATA_TEMPR56[1] ), .B(\R_DATA_TEMPR57[1] ), .C(
        \R_DATA_TEMPR58[1] ), .D(\R_DATA_TEMPR59[1] ), .Y(OR4_1188_Y));
    OR4 OR4_420 (.A(\R_DATA_TEMPR108[26] ), .B(\R_DATA_TEMPR109[26] ), 
        .C(\R_DATA_TEMPR110[26] ), .D(\R_DATA_TEMPR111[26] ), .Y(
        OR4_420_Y));
    OR4 OR4_738 (.A(OR4_1598_Y), .B(OR4_1438_Y), .C(OR4_1548_Y), .D(
        OR4_1149_Y), .Y(OR4_738_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[1]  (.A(CFG3_15_Y), .B(CFG3_2_Y)
        , .Y(\BLKY2[1] ));
    OR4 OR4_1141 (.A(\R_DATA_TEMPR40[18] ), .B(\R_DATA_TEMPR41[18] ), 
        .C(\R_DATA_TEMPR42[18] ), .D(\R_DATA_TEMPR43[18] ), .Y(
        OR4_1141_Y));
    OR4 OR4_402 (.A(\R_DATA_TEMPR116[36] ), .B(\R_DATA_TEMPR117[36] ), 
        .C(\R_DATA_TEMPR118[36] ), .D(\R_DATA_TEMPR119[36] ), .Y(
        OR4_402_Y));
    OR4 OR4_384 (.A(\R_DATA_TEMPR8[37] ), .B(\R_DATA_TEMPR9[37] ), .C(
        \R_DATA_TEMPR10[37] ), .D(\R_DATA_TEMPR11[37] ), .Y(OR4_384_Y));
    OR4 OR4_373 (.A(\R_DATA_TEMPR88[27] ), .B(\R_DATA_TEMPR89[27] ), 
        .C(\R_DATA_TEMPR90[27] ), .D(\R_DATA_TEMPR91[27] ), .Y(
        OR4_373_Y));
    OR4 OR4_770 (.A(\R_DATA_TEMPR116[16] ), .B(\R_DATA_TEMPR117[16] ), 
        .C(\R_DATA_TEMPR118[16] ), .D(\R_DATA_TEMPR119[16] ), .Y(
        OR4_770_Y));
    OR4 OR4_253 (.A(\R_DATA_TEMPR100[21] ), .B(\R_DATA_TEMPR101[21] ), 
        .C(\R_DATA_TEMPR102[21] ), .D(\R_DATA_TEMPR103[21] ), .Y(
        OR4_253_Y));
    OR4 OR4_1331 (.A(OR4_1502_Y), .B(OR4_23_Y), .C(OR4_143_Y), .D(
        OR4_33_Y), .Y(OR4_1331_Y));
    OR4 OR4_1463 (.A(OR4_697_Y), .B(OR4_149_Y), .C(OR4_122_Y), .D(
        OR4_912_Y), .Y(OR4_1463_Y));
    OR4 OR4_1253 (.A(\R_DATA_TEMPR96[2] ), .B(\R_DATA_TEMPR97[2] ), .C(
        \R_DATA_TEMPR98[2] ), .D(\R_DATA_TEMPR99[2] ), .Y(OR4_1253_Y));
    OR4 OR4_409 (.A(\R_DATA_TEMPR100[14] ), .B(\R_DATA_TEMPR101[14] ), 
        .C(\R_DATA_TEMPR102[14] ), .D(\R_DATA_TEMPR103[14] ), .Y(
        OR4_409_Y));
    OR4 OR4_472 (.A(\R_DATA_TEMPR0[1] ), .B(\R_DATA_TEMPR1[1] ), .C(
        \R_DATA_TEMPR2[1] ), .D(\R_DATA_TEMPR3[1] ), .Y(OR4_472_Y));
    OR4 OR4_1546 (.A(\R_DATA_TEMPR68[17] ), .B(\R_DATA_TEMPR69[17] ), 
        .C(\R_DATA_TEMPR70[17] ), .D(\R_DATA_TEMPR71[17] ), .Y(
        OR4_1546_Y));
    OR4 OR4_181 (.A(OR4_1179_Y), .B(OR4_1003_Y), .C(OR4_413_Y), .D(
        OR4_920_Y), .Y(OR4_181_Y));
    OR4 OR4_961 (.A(\R_DATA_TEMPR48[8] ), .B(\R_DATA_TEMPR49[8] ), .C(
        \R_DATA_TEMPR50[8] ), .D(\R_DATA_TEMPR51[8] ), .Y(OR4_961_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%64%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R64C0 (.A_DOUT({
        \R_DATA_TEMPR64[39] , \R_DATA_TEMPR64[38] , 
        \R_DATA_TEMPR64[37] , \R_DATA_TEMPR64[36] , 
        \R_DATA_TEMPR64[35] , \R_DATA_TEMPR64[34] , 
        \R_DATA_TEMPR64[33] , \R_DATA_TEMPR64[32] , 
        \R_DATA_TEMPR64[31] , \R_DATA_TEMPR64[30] , 
        \R_DATA_TEMPR64[29] , \R_DATA_TEMPR64[28] , 
        \R_DATA_TEMPR64[27] , \R_DATA_TEMPR64[26] , 
        \R_DATA_TEMPR64[25] , \R_DATA_TEMPR64[24] , 
        \R_DATA_TEMPR64[23] , \R_DATA_TEMPR64[22] , 
        \R_DATA_TEMPR64[21] , \R_DATA_TEMPR64[20] }), .B_DOUT({
        \R_DATA_TEMPR64[19] , \R_DATA_TEMPR64[18] , 
        \R_DATA_TEMPR64[17] , \R_DATA_TEMPR64[16] , 
        \R_DATA_TEMPR64[15] , \R_DATA_TEMPR64[14] , 
        \R_DATA_TEMPR64[13] , \R_DATA_TEMPR64[12] , 
        \R_DATA_TEMPR64[11] , \R_DATA_TEMPR64[10] , 
        \R_DATA_TEMPR64[9] , \R_DATA_TEMPR64[8] , \R_DATA_TEMPR64[7] , 
        \R_DATA_TEMPR64[6] , \R_DATA_TEMPR64[5] , \R_DATA_TEMPR64[4] , 
        \R_DATA_TEMPR64[3] , \R_DATA_TEMPR64[2] , \R_DATA_TEMPR64[1] , 
        \R_DATA_TEMPR64[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[64][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[16] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[16] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_106 (.A(\R_DATA_TEMPR0[6] ), .B(\R_DATA_TEMPR1[6] ), .C(
        \R_DATA_TEMPR2[6] ), .D(\R_DATA_TEMPR3[6] ), .Y(OR4_106_Y));
    OR4 OR4_958 (.A(\R_DATA_TEMPR80[30] ), .B(\R_DATA_TEMPR81[30] ), 
        .C(\R_DATA_TEMPR82[30] ), .D(\R_DATA_TEMPR83[30] ), .Y(
        OR4_958_Y));
    OR4 OR4_83 (.A(\R_DATA_TEMPR64[31] ), .B(\R_DATA_TEMPR65[31] ), .C(
        \R_DATA_TEMPR66[31] ), .D(\R_DATA_TEMPR67[31] ), .Y(OR4_83_Y));
    OR4 OR4_479 (.A(OR4_760_Y), .B(OR4_600_Y), .C(OR4_719_Y), .D(
        OR4_1419_Y), .Y(OR4_479_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[22]  (.A(CFG3_10_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[22] ));
    OR4 OR4_837 (.A(\R_DATA_TEMPR80[37] ), .B(\R_DATA_TEMPR81[37] ), 
        .C(\R_DATA_TEMPR82[37] ), .D(\R_DATA_TEMPR83[37] ), .Y(
        OR4_837_Y));
    OR4 OR4_138 (.A(\R_DATA_TEMPR68[14] ), .B(\R_DATA_TEMPR69[14] ), 
        .C(\R_DATA_TEMPR70[14] ), .D(\R_DATA_TEMPR71[14] ), .Y(
        OR4_138_Y));
    OR4 OR4_934 (.A(\R_DATA_TEMPR56[27] ), .B(\R_DATA_TEMPR57[27] ), 
        .C(\R_DATA_TEMPR58[27] ), .D(\R_DATA_TEMPR59[27] ), .Y(
        OR4_934_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%28%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C0 (.A_DOUT({
        \R_DATA_TEMPR28[39] , \R_DATA_TEMPR28[38] , 
        \R_DATA_TEMPR28[37] , \R_DATA_TEMPR28[36] , 
        \R_DATA_TEMPR28[35] , \R_DATA_TEMPR28[34] , 
        \R_DATA_TEMPR28[33] , \R_DATA_TEMPR28[32] , 
        \R_DATA_TEMPR28[31] , \R_DATA_TEMPR28[30] , 
        \R_DATA_TEMPR28[29] , \R_DATA_TEMPR28[28] , 
        \R_DATA_TEMPR28[27] , \R_DATA_TEMPR28[26] , 
        \R_DATA_TEMPR28[25] , \R_DATA_TEMPR28[24] , 
        \R_DATA_TEMPR28[23] , \R_DATA_TEMPR28[22] , 
        \R_DATA_TEMPR28[21] , \R_DATA_TEMPR28[20] }), .B_DOUT({
        \R_DATA_TEMPR28[19] , \R_DATA_TEMPR28[18] , 
        \R_DATA_TEMPR28[17] , \R_DATA_TEMPR28[16] , 
        \R_DATA_TEMPR28[15] , \R_DATA_TEMPR28[14] , 
        \R_DATA_TEMPR28[13] , \R_DATA_TEMPR28[12] , 
        \R_DATA_TEMPR28[11] , \R_DATA_TEMPR28[10] , 
        \R_DATA_TEMPR28[9] , \R_DATA_TEMPR28[8] , \R_DATA_TEMPR28[7] , 
        \R_DATA_TEMPR28[6] , \R_DATA_TEMPR28[5] , \R_DATA_TEMPR28[4] , 
        \R_DATA_TEMPR28[3] , \R_DATA_TEMPR28[2] , \R_DATA_TEMPR28[1] , 
        \R_DATA_TEMPR28[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1515 (.A(\R_DATA_TEMPR28[24] ), .B(\R_DATA_TEMPR29[24] ), 
        .C(\R_DATA_TEMPR30[24] ), .D(\R_DATA_TEMPR31[24] ), .Y(
        OR4_1515_Y));
    OR4 OR4_176 (.A(OR4_1109_Y), .B(OR4_735_Y), .C(OR4_704_Y), .D(
        OR4_1498_Y), .Y(OR4_176_Y));
    OR4 OR4_610 (.A(\R_DATA_TEMPR40[19] ), .B(\R_DATA_TEMPR41[19] ), 
        .C(\R_DATA_TEMPR42[19] ), .D(\R_DATA_TEMPR43[19] ), .Y(
        OR4_610_Y));
    OR4 OR4_481 (.A(\R_DATA_TEMPR120[17] ), .B(\R_DATA_TEMPR121[17] ), 
        .C(\R_DATA_TEMPR122[17] ), .D(\R_DATA_TEMPR123[17] ), .Y(
        OR4_481_Y));
    OR4 OR4_1216 (.A(\R_DATA_TEMPR96[24] ), .B(\R_DATA_TEMPR97[24] ), 
        .C(\R_DATA_TEMPR98[24] ), .D(\R_DATA_TEMPR99[24] ), .Y(
        OR4_1216_Y));
    OR4 OR4_1447 (.A(\R_DATA_TEMPR68[22] ), .B(\R_DATA_TEMPR69[22] ), 
        .C(\R_DATA_TEMPR70[22] ), .D(\R_DATA_TEMPR71[22] ), .Y(
        OR4_1447_Y));
    OR4 OR4_488 (.A(\R_DATA_TEMPR0[38] ), .B(\R_DATA_TEMPR1[38] ), .C(
        \R_DATA_TEMPR2[38] ), .D(\R_DATA_TEMPR3[38] ), .Y(OR4_488_Y));
    OR4 OR4_1072 (.A(\R_DATA_TEMPR56[29] ), .B(\R_DATA_TEMPR57[29] ), 
        .C(\R_DATA_TEMPR58[29] ), .D(\R_DATA_TEMPR59[29] ), .Y(
        OR4_1072_Y));
    OR4 OR4_308 (.A(OR4_749_Y), .B(OR2_38_Y), .C(\R_DATA_TEMPR86[10] ), 
        .D(\R_DATA_TEMPR87[10] ), .Y(OR4_308_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%117%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R117C0 (.A_DOUT({
        \R_DATA_TEMPR117[39] , \R_DATA_TEMPR117[38] , 
        \R_DATA_TEMPR117[37] , \R_DATA_TEMPR117[36] , 
        \R_DATA_TEMPR117[35] , \R_DATA_TEMPR117[34] , 
        \R_DATA_TEMPR117[33] , \R_DATA_TEMPR117[32] , 
        \R_DATA_TEMPR117[31] , \R_DATA_TEMPR117[30] , 
        \R_DATA_TEMPR117[29] , \R_DATA_TEMPR117[28] , 
        \R_DATA_TEMPR117[27] , \R_DATA_TEMPR117[26] , 
        \R_DATA_TEMPR117[25] , \R_DATA_TEMPR117[24] , 
        \R_DATA_TEMPR117[23] , \R_DATA_TEMPR117[22] , 
        \R_DATA_TEMPR117[21] , \R_DATA_TEMPR117[20] }), .B_DOUT({
        \R_DATA_TEMPR117[19] , \R_DATA_TEMPR117[18] , 
        \R_DATA_TEMPR117[17] , \R_DATA_TEMPR117[16] , 
        \R_DATA_TEMPR117[15] , \R_DATA_TEMPR117[14] , 
        \R_DATA_TEMPR117[13] , \R_DATA_TEMPR117[12] , 
        \R_DATA_TEMPR117[11] , \R_DATA_TEMPR117[10] , 
        \R_DATA_TEMPR117[9] , \R_DATA_TEMPR117[8] , 
        \R_DATA_TEMPR117[7] , \R_DATA_TEMPR117[6] , 
        \R_DATA_TEMPR117[5] , \R_DATA_TEMPR117[4] , 
        \R_DATA_TEMPR117[3] , \R_DATA_TEMPR117[2] , 
        \R_DATA_TEMPR117[1] , \R_DATA_TEMPR117[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[117][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[29] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[29] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1159 (.A(\R_DATA_TEMPR8[2] ), .B(\R_DATA_TEMPR9[2] ), .C(
        \R_DATA_TEMPR10[2] ), .D(\R_DATA_TEMPR11[2] ), .Y(OR4_1159_Y));
    OR4 OR4_317 (.A(\R_DATA_TEMPR56[22] ), .B(\R_DATA_TEMPR57[22] ), 
        .C(\R_DATA_TEMPR58[22] ), .D(\R_DATA_TEMPR59[22] ), .Y(
        OR4_317_Y));
    OR4 OR4_110 (.A(\R_DATA_TEMPR88[12] ), .B(\R_DATA_TEMPR89[12] ), 
        .C(\R_DATA_TEMPR90[12] ), .D(\R_DATA_TEMPR91[12] ), .Y(
        OR4_110_Y));
    OR4 OR4_848 (.A(\R_DATA_TEMPR36[39] ), .B(\R_DATA_TEMPR37[39] ), 
        .C(\R_DATA_TEMPR38[39] ), .D(\R_DATA_TEMPR39[39] ), .Y(
        OR4_848_Y));
    OR4 OR4_1318 (.A(\R_DATA_TEMPR36[33] ), .B(\R_DATA_TEMPR37[33] ), 
        .C(\R_DATA_TEMPR38[33] ), .D(\R_DATA_TEMPR39[33] ), .Y(
        OR4_1318_Y));
    CFG3 #( .INIT(8'h1) )  CFG3_16 (.A(R_ADDR[13]), .B(R_ADDR[12]), .C(
        R_ADDR[11]), .Y(CFG3_16_Y));
    OR4 OR4_1026 (.A(OR4_840_Y), .B(OR2_7_Y), .C(\R_DATA_TEMPR86[28] ), 
        .D(\R_DATA_TEMPR87[28] ), .Y(OR4_1026_Y));
    OR4 OR4_658 (.A(\R_DATA_TEMPR64[4] ), .B(\R_DATA_TEMPR65[4] ), .C(
        \R_DATA_TEMPR66[4] ), .D(\R_DATA_TEMPR67[4] ), .Y(OR4_658_Y));
    OR4 OR4_1045 (.A(OR4_811_Y), .B(OR4_1632_Y), .C(OR4_540_Y), .D(
        OR4_1564_Y), .Y(OR4_1045_Y));
    OR4 OR4_799 (.A(\R_DATA_TEMPR96[38] ), .B(\R_DATA_TEMPR97[38] ), 
        .C(\R_DATA_TEMPR98[38] ), .D(\R_DATA_TEMPR99[38] ), .Y(
        OR4_799_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%31%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C0 (.A_DOUT({
        \R_DATA_TEMPR31[39] , \R_DATA_TEMPR31[38] , 
        \R_DATA_TEMPR31[37] , \R_DATA_TEMPR31[36] , 
        \R_DATA_TEMPR31[35] , \R_DATA_TEMPR31[34] , 
        \R_DATA_TEMPR31[33] , \R_DATA_TEMPR31[32] , 
        \R_DATA_TEMPR31[31] , \R_DATA_TEMPR31[30] , 
        \R_DATA_TEMPR31[29] , \R_DATA_TEMPR31[28] , 
        \R_DATA_TEMPR31[27] , \R_DATA_TEMPR31[26] , 
        \R_DATA_TEMPR31[25] , \R_DATA_TEMPR31[24] , 
        \R_DATA_TEMPR31[23] , \R_DATA_TEMPR31[22] , 
        \R_DATA_TEMPR31[21] , \R_DATA_TEMPR31[20] }), .B_DOUT({
        \R_DATA_TEMPR31[19] , \R_DATA_TEMPR31[18] , 
        \R_DATA_TEMPR31[17] , \R_DATA_TEMPR31[16] , 
        \R_DATA_TEMPR31[15] , \R_DATA_TEMPR31[14] , 
        \R_DATA_TEMPR31[13] , \R_DATA_TEMPR31[12] , 
        \R_DATA_TEMPR31[11] , \R_DATA_TEMPR31[10] , 
        \R_DATA_TEMPR31[9] , \R_DATA_TEMPR31[8] , \R_DATA_TEMPR31[7] , 
        \R_DATA_TEMPR31[6] , \R_DATA_TEMPR31[5] , \R_DATA_TEMPR31[4] , 
        \R_DATA_TEMPR31[3] , \R_DATA_TEMPR31[2] , \R_DATA_TEMPR31[1] , 
        \R_DATA_TEMPR31[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_378 (.A(OR4_1083_Y), .B(OR4_1609_Y), .C(OR4_1107_Y), .D(
        OR4_612_Y), .Y(OR4_378_Y));
    OR4 OR4_2 (.A(OR4_568_Y), .B(OR4_835_Y), .C(OR4_828_Y), .D(
        OR4_1096_Y), .Y(OR4_2_Y));
    OR4 OR4_718 (.A(OR4_748_Y), .B(OR4_1051_Y), .C(OR4_513_Y), .D(
        OR4_1367_Y), .Y(OR4_718_Y));
    OR4 OR4_329 (.A(\R_DATA_TEMPR64[14] ), .B(\R_DATA_TEMPR65[14] ), 
        .C(\R_DATA_TEMPR66[14] ), .D(\R_DATA_TEMPR67[14] ), .Y(
        OR4_329_Y));
    OR4 \OR4_R_DATA[29]  (.A(OR4_390_Y), .B(OR4_20_Y), .C(OR4_1543_Y), 
        .D(OR4_1266_Y), .Y(R_DATA[29]));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%7%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C0 (.A_DOUT({
        \R_DATA_TEMPR7[39] , \R_DATA_TEMPR7[38] , \R_DATA_TEMPR7[37] , 
        \R_DATA_TEMPR7[36] , \R_DATA_TEMPR7[35] , \R_DATA_TEMPR7[34] , 
        \R_DATA_TEMPR7[33] , \R_DATA_TEMPR7[32] , \R_DATA_TEMPR7[31] , 
        \R_DATA_TEMPR7[30] , \R_DATA_TEMPR7[29] , \R_DATA_TEMPR7[28] , 
        \R_DATA_TEMPR7[27] , \R_DATA_TEMPR7[26] , \R_DATA_TEMPR7[25] , 
        \R_DATA_TEMPR7[24] , \R_DATA_TEMPR7[23] , \R_DATA_TEMPR7[22] , 
        \R_DATA_TEMPR7[21] , \R_DATA_TEMPR7[20] }), .B_DOUT({
        \R_DATA_TEMPR7[19] , \R_DATA_TEMPR7[18] , \R_DATA_TEMPR7[17] , 
        \R_DATA_TEMPR7[16] , \R_DATA_TEMPR7[15] , \R_DATA_TEMPR7[14] , 
        \R_DATA_TEMPR7[13] , \R_DATA_TEMPR7[12] , \R_DATA_TEMPR7[11] , 
        \R_DATA_TEMPR7[10] , \R_DATA_TEMPR7[9] , \R_DATA_TEMPR7[8] , 
        \R_DATA_TEMPR7[7] , \R_DATA_TEMPR7[6] , \R_DATA_TEMPR7[5] , 
        \R_DATA_TEMPR7[4] , \R_DATA_TEMPR7[3] , \R_DATA_TEMPR7[2] , 
        \R_DATA_TEMPR7[1] , \R_DATA_TEMPR7[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[7][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_894 (.A(\R_DATA_TEMPR112[36] ), .B(\R_DATA_TEMPR113[36] ), 
        .C(\R_DATA_TEMPR114[36] ), .D(\R_DATA_TEMPR115[36] ), .Y(
        OR4_894_Y));
    OR4 OR4_765 (.A(\R_DATA_TEMPR48[18] ), .B(\R_DATA_TEMPR49[18] ), 
        .C(\R_DATA_TEMPR50[18] ), .D(\R_DATA_TEMPR51[18] ), .Y(
        OR4_765_Y));
    OR4 OR4_667 (.A(\R_DATA_TEMPR16[35] ), .B(\R_DATA_TEMPR17[35] ), 
        .C(\R_DATA_TEMPR18[35] ), .D(\R_DATA_TEMPR19[35] ), .Y(
        OR4_667_Y));
    OR4 OR4_652 (.A(\R_DATA_TEMPR16[11] ), .B(\R_DATA_TEMPR17[11] ), 
        .C(\R_DATA_TEMPR18[11] ), .D(\R_DATA_TEMPR19[11] ), .Y(
        OR4_652_Y));
    OR4 OR4_1493 (.A(\R_DATA_TEMPR100[13] ), .B(\R_DATA_TEMPR101[13] ), 
        .C(\R_DATA_TEMPR102[13] ), .D(\R_DATA_TEMPR103[13] ), .Y(
        OR4_1493_Y));
    OR4 OR4_1321 (.A(\R_DATA_TEMPR112[29] ), .B(\R_DATA_TEMPR113[29] ), 
        .C(\R_DATA_TEMPR114[29] ), .D(\R_DATA_TEMPR115[29] ), .Y(
        OR4_1321_Y));
    OR4 OR4_766 (.A(OR4_1549_Y), .B(OR4_1058_Y), .C(OR4_1139_Y), .D(
        OR4_1456_Y), .Y(OR4_766_Y));
    OR4 OR4_593 (.A(\R_DATA_TEMPR108[4] ), .B(\R_DATA_TEMPR109[4] ), 
        .C(\R_DATA_TEMPR110[4] ), .D(\R_DATA_TEMPR111[4] ), .Y(
        OR4_593_Y));
    OR4 OR4_48 (.A(\R_DATA_TEMPR120[14] ), .B(\R_DATA_TEMPR121[14] ), 
        .C(\R_DATA_TEMPR122[14] ), .D(\R_DATA_TEMPR123[14] ), .Y(
        OR4_48_Y));
    OR4 OR4_589 (.A(OR4_1516_Y), .B(OR2_28_Y), .C(\R_DATA_TEMPR86[35] )
        , .D(\R_DATA_TEMPR87[35] ), .Y(OR4_589_Y));
    OR2 OR2_33 (.A(\R_DATA_TEMPR84[6] ), .B(\R_DATA_TEMPR85[6] ), .Y(
        OR2_33_Y));
    OR4 OR4_109 (.A(\R_DATA_TEMPR52[1] ), .B(\R_DATA_TEMPR53[1] ), .C(
        \R_DATA_TEMPR54[1] ), .D(\R_DATA_TEMPR55[1] ), .Y(OR4_109_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%94%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R94C0 (.A_DOUT({
        \R_DATA_TEMPR94[39] , \R_DATA_TEMPR94[38] , 
        \R_DATA_TEMPR94[37] , \R_DATA_TEMPR94[36] , 
        \R_DATA_TEMPR94[35] , \R_DATA_TEMPR94[34] , 
        \R_DATA_TEMPR94[33] , \R_DATA_TEMPR94[32] , 
        \R_DATA_TEMPR94[31] , \R_DATA_TEMPR94[30] , 
        \R_DATA_TEMPR94[29] , \R_DATA_TEMPR94[28] , 
        \R_DATA_TEMPR94[27] , \R_DATA_TEMPR94[26] , 
        \R_DATA_TEMPR94[25] , \R_DATA_TEMPR94[24] , 
        \R_DATA_TEMPR94[23] , \R_DATA_TEMPR94[22] , 
        \R_DATA_TEMPR94[21] , \R_DATA_TEMPR94[20] }), .B_DOUT({
        \R_DATA_TEMPR94[19] , \R_DATA_TEMPR94[18] , 
        \R_DATA_TEMPR94[17] , \R_DATA_TEMPR94[16] , 
        \R_DATA_TEMPR94[15] , \R_DATA_TEMPR94[14] , 
        \R_DATA_TEMPR94[13] , \R_DATA_TEMPR94[12] , 
        \R_DATA_TEMPR94[11] , \R_DATA_TEMPR94[10] , 
        \R_DATA_TEMPR94[9] , \R_DATA_TEMPR94[8] , \R_DATA_TEMPR94[7] , 
        \R_DATA_TEMPR94[6] , \R_DATA_TEMPR94[5] , \R_DATA_TEMPR94[4] , 
        \R_DATA_TEMPR94[3] , \R_DATA_TEMPR94[2] , \R_DATA_TEMPR94[1] , 
        \R_DATA_TEMPR94[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[94][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[23] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[23] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_15 (.A(\R_DATA_TEMPR84[8] ), .B(\R_DATA_TEMPR85[8] ), .Y(
        OR2_15_Y));
    OR4 OR4_241 (.A(\R_DATA_TEMPR20[18] ), .B(\R_DATA_TEMPR21[18] ), 
        .C(\R_DATA_TEMPR22[18] ), .D(\R_DATA_TEMPR23[18] ), .Y(
        OR4_241_Y));
    OR4 OR4_580 (.A(\R_DATA_TEMPR12[0] ), .B(\R_DATA_TEMPR13[0] ), .C(
        \R_DATA_TEMPR14[0] ), .D(\R_DATA_TEMPR15[0] ), .Y(OR4_580_Y));
    OR4 OR4_81 (.A(\R_DATA_TEMPR28[10] ), .B(\R_DATA_TEMPR29[10] ), .C(
        \R_DATA_TEMPR30[10] ), .D(\R_DATA_TEMPR31[10] ), .Y(OR4_81_Y));
    OR4 OR4_1019 (.A(\R_DATA_TEMPR48[34] ), .B(\R_DATA_TEMPR49[34] ), 
        .C(\R_DATA_TEMPR50[34] ), .D(\R_DATA_TEMPR51[34] ), .Y(
        OR4_1019_Y));
    OR4 OR4_817 (.A(\R_DATA_TEMPR68[10] ), .B(\R_DATA_TEMPR69[10] ), 
        .C(\R_DATA_TEMPR70[10] ), .D(\R_DATA_TEMPR71[10] ), .Y(
        OR4_817_Y));
    OR4 OR4_118 (.A(\R_DATA_TEMPR20[37] ), .B(\R_DATA_TEMPR21[37] ), 
        .C(\R_DATA_TEMPR22[37] ), .D(\R_DATA_TEMPR23[37] ), .Y(
        OR4_118_Y));
    OR4 OR4_914 (.A(\R_DATA_TEMPR56[30] ), .B(\R_DATA_TEMPR57[30] ), 
        .C(\R_DATA_TEMPR58[30] ), .D(\R_DATA_TEMPR59[30] ), .Y(
        OR4_914_Y));
    OR4 \OR4_R_DATA[7]  (.A(OR4_953_Y), .B(OR4_1499_Y), .C(OR4_1032_Y), 
        .D(OR4_800_Y), .Y(R_DATA[7]));
    OR4 OR4_179 (.A(\R_DATA_TEMPR20[3] ), .B(\R_DATA_TEMPR21[3] ), .C(
        \R_DATA_TEMPR22[3] ), .D(\R_DATA_TEMPR23[3] ), .Y(OR4_179_Y));
    OR4 OR4_1163 (.A(\R_DATA_TEMPR64[5] ), .B(\R_DATA_TEMPR65[5] ), .C(
        \R_DATA_TEMPR66[5] ), .D(\R_DATA_TEMPR67[5] ), .Y(OR4_1163_Y));
    OR4 OR4_1156 (.A(OR4_1490_Y), .B(OR4_848_Y), .C(OR4_823_Y), .D(
        OR4_514_Y), .Y(OR4_1156_Y));
    OR4 OR4_1451 (.A(\R_DATA_TEMPR104[1] ), .B(\R_DATA_TEMPR105[1] ), 
        .C(\R_DATA_TEMPR106[1] ), .D(\R_DATA_TEMPR107[1] ), .Y(
        OR4_1451_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%60%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R60C0 (.A_DOUT({
        \R_DATA_TEMPR60[39] , \R_DATA_TEMPR60[38] , 
        \R_DATA_TEMPR60[37] , \R_DATA_TEMPR60[36] , 
        \R_DATA_TEMPR60[35] , \R_DATA_TEMPR60[34] , 
        \R_DATA_TEMPR60[33] , \R_DATA_TEMPR60[32] , 
        \R_DATA_TEMPR60[31] , \R_DATA_TEMPR60[30] , 
        \R_DATA_TEMPR60[29] , \R_DATA_TEMPR60[28] , 
        \R_DATA_TEMPR60[27] , \R_DATA_TEMPR60[26] , 
        \R_DATA_TEMPR60[25] , \R_DATA_TEMPR60[24] , 
        \R_DATA_TEMPR60[23] , \R_DATA_TEMPR60[22] , 
        \R_DATA_TEMPR60[21] , \R_DATA_TEMPR60[20] }), .B_DOUT({
        \R_DATA_TEMPR60[19] , \R_DATA_TEMPR60[18] , 
        \R_DATA_TEMPR60[17] , \R_DATA_TEMPR60[16] , 
        \R_DATA_TEMPR60[15] , \R_DATA_TEMPR60[14] , 
        \R_DATA_TEMPR60[13] , \R_DATA_TEMPR60[12] , 
        \R_DATA_TEMPR60[11] , \R_DATA_TEMPR60[10] , 
        \R_DATA_TEMPR60[9] , \R_DATA_TEMPR60[8] , \R_DATA_TEMPR60[7] , 
        \R_DATA_TEMPR60[6] , \R_DATA_TEMPR60[5] , \R_DATA_TEMPR60[4] , 
        \R_DATA_TEMPR60[3] , \R_DATA_TEMPR60[2] , \R_DATA_TEMPR60[1] , 
        \R_DATA_TEMPR60[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[60][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[15] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[15] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1251 (.A(\R_DATA_TEMPR48[21] ), .B(\R_DATA_TEMPR49[21] ), 
        .C(\R_DATA_TEMPR50[21] ), .D(\R_DATA_TEMPR51[21] ), .Y(
        OR4_1251_Y));
    OR4 OR4_901 (.A(\R_DATA_TEMPR32[4] ), .B(\R_DATA_TEMPR33[4] ), .C(
        \R_DATA_TEMPR34[4] ), .D(\R_DATA_TEMPR35[4] ), .Y(OR4_901_Y));
    OR4 OR4_1158 (.A(\R_DATA_TEMPR112[13] ), .B(\R_DATA_TEMPR113[13] ), 
        .C(\R_DATA_TEMPR114[13] ), .D(\R_DATA_TEMPR115[13] ), .Y(
        OR4_1158_Y));
    OR4 OR4_542 (.A(\R_DATA_TEMPR68[32] ), .B(\R_DATA_TEMPR69[32] ), 
        .C(\R_DATA_TEMPR70[32] ), .D(\R_DATA_TEMPR71[32] ), .Y(
        OR4_542_Y));
    OR4 OR4_1132 (.A(OR4_837_Y), .B(OR2_12_Y), .C(\R_DATA_TEMPR86[37] )
        , .D(\R_DATA_TEMPR87[37] ), .Y(OR4_1132_Y));
    OR4 OR4_1569 (.A(OR4_431_Y), .B(OR4_885_Y), .C(OR4_217_Y), .D(
        OR4_532_Y), .Y(OR4_1569_Y));
    OR4 OR4_855 (.A(OR4_716_Y), .B(OR4_222_Y), .C(OR4_276_Y), .D(
        OR4_1618_Y), .Y(OR4_855_Y));
    OR4 OR4_971 (.A(OR4_1210_Y), .B(OR4_1485_Y), .C(OR4_17_Y), .D(
        OR4_903_Y), .Y(OR4_971_Y));
    OR4 OR4_1603 (.A(OR4_1404_Y), .B(OR4_1617_Y), .C(OR4_1596_Y), .D(
        OR4_1270_Y), .Y(OR4_1603_Y));
    OR4 OR4_1573 (.A(\R_DATA_TEMPR76[23] ), .B(\R_DATA_TEMPR77[23] ), 
        .C(\R_DATA_TEMPR78[23] ), .D(\R_DATA_TEMPR79[23] ), .Y(
        OR4_1573_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%27%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C0 (.A_DOUT({
        \R_DATA_TEMPR27[39] , \R_DATA_TEMPR27[38] , 
        \R_DATA_TEMPR27[37] , \R_DATA_TEMPR27[36] , 
        \R_DATA_TEMPR27[35] , \R_DATA_TEMPR27[34] , 
        \R_DATA_TEMPR27[33] , \R_DATA_TEMPR27[32] , 
        \R_DATA_TEMPR27[31] , \R_DATA_TEMPR27[30] , 
        \R_DATA_TEMPR27[29] , \R_DATA_TEMPR27[28] , 
        \R_DATA_TEMPR27[27] , \R_DATA_TEMPR27[26] , 
        \R_DATA_TEMPR27[25] , \R_DATA_TEMPR27[24] , 
        \R_DATA_TEMPR27[23] , \R_DATA_TEMPR27[22] , 
        \R_DATA_TEMPR27[21] , \R_DATA_TEMPR27[20] }), .B_DOUT({
        \R_DATA_TEMPR27[19] , \R_DATA_TEMPR27[18] , 
        \R_DATA_TEMPR27[17] , \R_DATA_TEMPR27[16] , 
        \R_DATA_TEMPR27[15] , \R_DATA_TEMPR27[14] , 
        \R_DATA_TEMPR27[13] , \R_DATA_TEMPR27[12] , 
        \R_DATA_TEMPR27[11] , \R_DATA_TEMPR27[10] , 
        \R_DATA_TEMPR27[9] , \R_DATA_TEMPR27[8] , \R_DATA_TEMPR27[7] , 
        \R_DATA_TEMPR27[6] , \R_DATA_TEMPR27[5] , \R_DATA_TEMPR27[4] , 
        \R_DATA_TEMPR27[3] , \R_DATA_TEMPR27[2] , \R_DATA_TEMPR27[1] , 
        \R_DATA_TEMPR27[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_729 (.A(\R_DATA_TEMPR104[20] ), .B(\R_DATA_TEMPR105[20] ), 
        .C(\R_DATA_TEMPR106[20] ), .D(\R_DATA_TEMPR107[20] ), .Y(
        OR4_729_Y));
    OR4 OR4_1504 (.A(\R_DATA_TEMPR76[26] ), .B(\R_DATA_TEMPR77[26] ), 
        .C(\R_DATA_TEMPR78[26] ), .D(\R_DATA_TEMPR79[26] ), .Y(
        OR4_1504_Y));
    OR4 \OR4_R_DATA[4]  (.A(OR4_1252_Y), .B(OR4_330_Y), .C(OR4_534_Y), 
        .D(OR4_707_Y), .Y(R_DATA[4]));
    OR4 OR4_135 (.A(OR4_97_Y), .B(OR4_409_Y), .C(OR4_647_Y), .D(
        OR4_461_Y), .Y(OR4_135_Y));
    OR4 OR4_824 (.A(\R_DATA_TEMPR20[7] ), .B(\R_DATA_TEMPR21[7] ), .C(
        \R_DATA_TEMPR22[7] ), .D(\R_DATA_TEMPR23[7] ), .Y(OR4_824_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[9]  (.A(CFG3_15_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[9] ));
    OR4 OR4_383 (.A(OR4_1309_Y), .B(OR2_10_Y), .C(\R_DATA_TEMPR86[15] )
        , .D(\R_DATA_TEMPR87[15] ), .Y(OR4_383_Y));
    OR4 OR4_1305 (.A(\R_DATA_TEMPR72[3] ), .B(\R_DATA_TEMPR73[3] ), .C(
        \R_DATA_TEMPR74[3] ), .D(\R_DATA_TEMPR75[3] ), .Y(OR4_1305_Y));
    OR4 OR4_1140 (.A(\R_DATA_TEMPR24[14] ), .B(\R_DATA_TEMPR25[14] ), 
        .C(\R_DATA_TEMPR26[14] ), .D(\R_DATA_TEMPR27[14] ), .Y(
        OR4_1140_Y));
    OR4 OR4_780 (.A(\R_DATA_TEMPR88[31] ), .B(\R_DATA_TEMPR89[31] ), 
        .C(\R_DATA_TEMPR90[31] ), .D(\R_DATA_TEMPR91[31] ), .Y(
        OR4_780_Y));
    OR4 OR4_544 (.A(OR4_1250_Y), .B(OR4_1327_Y), .C(OR4_1295_Y), .D(
        OR4_972_Y), .Y(OR4_544_Y));
    OR2 OR2_31 (.A(\R_DATA_TEMPR84[38] ), .B(\R_DATA_TEMPR85[38] ), .Y(
        OR2_31_Y));
    OR4 OR4_267 (.A(OR4_1163_Y), .B(OR4_1443_Y), .C(OR4_1628_Y), .D(
        OR4_1401_Y), .Y(OR4_267_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%4%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C0 (.A_DOUT({
        \R_DATA_TEMPR4[39] , \R_DATA_TEMPR4[38] , \R_DATA_TEMPR4[37] , 
        \R_DATA_TEMPR4[36] , \R_DATA_TEMPR4[35] , \R_DATA_TEMPR4[34] , 
        \R_DATA_TEMPR4[33] , \R_DATA_TEMPR4[32] , \R_DATA_TEMPR4[31] , 
        \R_DATA_TEMPR4[30] , \R_DATA_TEMPR4[29] , \R_DATA_TEMPR4[28] , 
        \R_DATA_TEMPR4[27] , \R_DATA_TEMPR4[26] , \R_DATA_TEMPR4[25] , 
        \R_DATA_TEMPR4[24] , \R_DATA_TEMPR4[23] , \R_DATA_TEMPR4[22] , 
        \R_DATA_TEMPR4[21] , \R_DATA_TEMPR4[20] }), .B_DOUT({
        \R_DATA_TEMPR4[19] , \R_DATA_TEMPR4[18] , \R_DATA_TEMPR4[17] , 
        \R_DATA_TEMPR4[16] , \R_DATA_TEMPR4[15] , \R_DATA_TEMPR4[14] , 
        \R_DATA_TEMPR4[13] , \R_DATA_TEMPR4[12] , \R_DATA_TEMPR4[11] , 
        \R_DATA_TEMPR4[10] , \R_DATA_TEMPR4[9] , \R_DATA_TEMPR4[8] , 
        \R_DATA_TEMPR4[7] , \R_DATA_TEMPR4[6] , \R_DATA_TEMPR4[5] , 
        \R_DATA_TEMPR4[4] , \R_DATA_TEMPR4[3] , \R_DATA_TEMPR4[2] , 
        \R_DATA_TEMPR4[1] , \R_DATA_TEMPR4[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[4][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h8) )  CFG3_9 (.A(R_EN), .B(R_ADDR[15]), .C(
        R_ADDR[14]), .Y(CFG3_9_Y));
    OR4 OR4_523 (.A(\R_DATA_TEMPR112[6] ), .B(\R_DATA_TEMPR113[6] ), 
        .C(\R_DATA_TEMPR114[6] ), .D(\R_DATA_TEMPR115[6] ), .Y(
        OR4_523_Y));
    OR4 OR4_437 (.A(\R_DATA_TEMPR44[5] ), .B(\R_DATA_TEMPR45[5] ), .C(
        \R_DATA_TEMPR46[5] ), .D(\R_DATA_TEMPR47[5] ), .Y(OR4_437_Y));
    OR4 OR4_942 (.A(\R_DATA_TEMPR4[5] ), .B(\R_DATA_TEMPR5[5] ), .C(
        \R_DATA_TEMPR6[5] ), .D(\R_DATA_TEMPR7[5] ), .Y(OR4_942_Y));
    OR4 OR4_482 (.A(\R_DATA_TEMPR48[16] ), .B(\R_DATA_TEMPR49[16] ), 
        .C(\R_DATA_TEMPR50[16] ), .D(\R_DATA_TEMPR51[16] ), .Y(
        OR4_482_Y));
    OR4 OR4_167 (.A(\R_DATA_TEMPR56[6] ), .B(\R_DATA_TEMPR57[6] ), .C(
        \R_DATA_TEMPR58[6] ), .D(\R_DATA_TEMPR59[6] ), .Y(OR4_167_Y));
    OR4 OR4_1193 (.A(OR4_444_Y), .B(OR4_1079_Y), .C(OR4_1620_Y), .D(
        OR4_439_Y), .Y(OR4_1193_Y));
    OR4 OR4_705 (.A(\R_DATA_TEMPR92[13] ), .B(\R_DATA_TEMPR93[13] ), 
        .C(\R_DATA_TEMPR94[13] ), .D(\R_DATA_TEMPR95[13] ), .Y(
        OR4_705_Y));
    OR4 OR4_607 (.A(\R_DATA_TEMPR124[16] ), .B(\R_DATA_TEMPR125[16] ), 
        .C(\R_DATA_TEMPR126[16] ), .D(\R_DATA_TEMPR127[16] ), .Y(
        OR4_607_Y));
    OR4 OR4_489 (.A(OR4_483_Y), .B(OR2_36_Y), .C(\R_DATA_TEMPR86[23] ), 
        .D(\R_DATA_TEMPR87[23] ), .Y(OR4_489_Y));
    OR4 OR4_706 (.A(\R_DATA_TEMPR28[4] ), .B(\R_DATA_TEMPR29[4] ), .C(
        \R_DATA_TEMPR30[4] ), .D(\R_DATA_TEMPR31[4] ), .Y(OR4_706_Y));
    OR4 OR4_186 (.A(OR4_1507_Y), .B(OR4_1344_Y), .C(OR4_1482_Y), .D(
        OR4_664_Y), .Y(OR4_186_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%90%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R90C0 (.A_DOUT({
        \R_DATA_TEMPR90[39] , \R_DATA_TEMPR90[38] , 
        \R_DATA_TEMPR90[37] , \R_DATA_TEMPR90[36] , 
        \R_DATA_TEMPR90[35] , \R_DATA_TEMPR90[34] , 
        \R_DATA_TEMPR90[33] , \R_DATA_TEMPR90[32] , 
        \R_DATA_TEMPR90[31] , \R_DATA_TEMPR90[30] , 
        \R_DATA_TEMPR90[29] , \R_DATA_TEMPR90[28] , 
        \R_DATA_TEMPR90[27] , \R_DATA_TEMPR90[26] , 
        \R_DATA_TEMPR90[25] , \R_DATA_TEMPR90[24] , 
        \R_DATA_TEMPR90[23] , \R_DATA_TEMPR90[22] , 
        \R_DATA_TEMPR90[21] , \R_DATA_TEMPR90[20] }), .B_DOUT({
        \R_DATA_TEMPR90[19] , \R_DATA_TEMPR90[18] , 
        \R_DATA_TEMPR90[17] , \R_DATA_TEMPR90[16] , 
        \R_DATA_TEMPR90[15] , \R_DATA_TEMPR90[14] , 
        \R_DATA_TEMPR90[13] , \R_DATA_TEMPR90[12] , 
        \R_DATA_TEMPR90[11] , \R_DATA_TEMPR90[10] , 
        \R_DATA_TEMPR90[9] , \R_DATA_TEMPR90[8] , \R_DATA_TEMPR90[7] , 
        \R_DATA_TEMPR90[6] , \R_DATA_TEMPR90[5] , \R_DATA_TEMPR90[4] , 
        \R_DATA_TEMPR90[3] , \R_DATA_TEMPR90[2] , \R_DATA_TEMPR90[1] , 
        \R_DATA_TEMPR90[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[90][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[22] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[22] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_775 (.A(\R_DATA_TEMPR116[6] ), .B(\R_DATA_TEMPR117[6] ), 
        .C(\R_DATA_TEMPR118[6] ), .D(\R_DATA_TEMPR119[6] ), .Y(
        OR4_775_Y));
    OR4 OR4_677 (.A(\R_DATA_TEMPR120[33] ), .B(\R_DATA_TEMPR121[33] ), 
        .C(\R_DATA_TEMPR122[33] ), .D(\R_DATA_TEMPR123[33] ), .Y(
        OR4_677_Y));
    OR4 OR4_1584 (.A(\R_DATA_TEMPR0[21] ), .B(\R_DATA_TEMPR1[21] ), .C(
        \R_DATA_TEMPR2[21] ), .D(\R_DATA_TEMPR3[21] ), .Y(OR4_1584_Y));
    OR4 OR4_235 (.A(\R_DATA_TEMPR8[25] ), .B(\R_DATA_TEMPR9[25] ), .C(
        \R_DATA_TEMPR10[25] ), .D(\R_DATA_TEMPR11[25] ), .Y(OR4_235_Y));
    OR4 OR4_341 (.A(\R_DATA_TEMPR40[26] ), .B(\R_DATA_TEMPR41[26] ), 
        .C(\R_DATA_TEMPR42[26] ), .D(\R_DATA_TEMPR43[26] ), .Y(
        OR4_341_Y));
    OR4 OR4_1599 (.A(\R_DATA_TEMPR124[5] ), .B(\R_DATA_TEMPR125[5] ), 
        .C(\R_DATA_TEMPR126[5] ), .D(\R_DATA_TEMPR127[5] ), .Y(
        OR4_1599_Y));
    OR4 OR4_776 (.A(\R_DATA_TEMPR56[19] ), .B(\R_DATA_TEMPR57[19] ), 
        .C(\R_DATA_TEMPR58[19] ), .D(\R_DATA_TEMPR59[19] ), .Y(
        OR4_776_Y));
    OR4 OR4_1122 (.A(\R_DATA_TEMPR0[15] ), .B(\R_DATA_TEMPR1[15] ), .C(
        \R_DATA_TEMPR2[15] ), .D(\R_DATA_TEMPR3[15] ), .Y(OR4_1122_Y));
    OR4 OR4_763 (.A(\R_DATA_TEMPR28[37] ), .B(\R_DATA_TEMPR29[37] ), 
        .C(\R_DATA_TEMPR30[37] ), .D(\R_DATA_TEMPR31[37] ), .Y(
        OR4_763_Y));
    OR2 OR2_29 (.A(\R_DATA_TEMPR84[22] ), .B(\R_DATA_TEMPR85[22] ), .Y(
        OR2_29_Y));
    OR4 OR4_832 (.A(\R_DATA_TEMPR108[22] ), .B(\R_DATA_TEMPR109[22] ), 
        .C(\R_DATA_TEMPR110[22] ), .D(\R_DATA_TEMPR111[22] ), .Y(
        OR4_832_Y));
    OR4 OR4_1565 (.A(\R_DATA_TEMPR28[11] ), .B(\R_DATA_TEMPR29[11] ), 
        .C(\R_DATA_TEMPR30[11] ), .D(\R_DATA_TEMPR31[11] ), .Y(
        OR4_1565_Y));
    OR4 OR4_1385 (.A(\R_DATA_TEMPR48[15] ), .B(\R_DATA_TEMPR49[15] ), 
        .C(\R_DATA_TEMPR50[15] ), .D(\R_DATA_TEMPR51[15] ), .Y(
        OR4_1385_Y));
    OR4 OR4_264 (.A(OR4_204_Y), .B(OR2_19_Y), .C(\R_DATA_TEMPR86[9] ), 
        .D(\R_DATA_TEMPR87[9] ), .Y(OR4_264_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%73%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R73C0 (.A_DOUT({
        \R_DATA_TEMPR73[39] , \R_DATA_TEMPR73[38] , 
        \R_DATA_TEMPR73[37] , \R_DATA_TEMPR73[36] , 
        \R_DATA_TEMPR73[35] , \R_DATA_TEMPR73[34] , 
        \R_DATA_TEMPR73[33] , \R_DATA_TEMPR73[32] , 
        \R_DATA_TEMPR73[31] , \R_DATA_TEMPR73[30] , 
        \R_DATA_TEMPR73[29] , \R_DATA_TEMPR73[28] , 
        \R_DATA_TEMPR73[27] , \R_DATA_TEMPR73[26] , 
        \R_DATA_TEMPR73[25] , \R_DATA_TEMPR73[24] , 
        \R_DATA_TEMPR73[23] , \R_DATA_TEMPR73[22] , 
        \R_DATA_TEMPR73[21] , \R_DATA_TEMPR73[20] }), .B_DOUT({
        \R_DATA_TEMPR73[19] , \R_DATA_TEMPR73[18] , 
        \R_DATA_TEMPR73[17] , \R_DATA_TEMPR73[16] , 
        \R_DATA_TEMPR73[15] , \R_DATA_TEMPR73[14] , 
        \R_DATA_TEMPR73[13] , \R_DATA_TEMPR73[12] , 
        \R_DATA_TEMPR73[11] , \R_DATA_TEMPR73[10] , 
        \R_DATA_TEMPR73[9] , \R_DATA_TEMPR73[8] , \R_DATA_TEMPR73[7] , 
        \R_DATA_TEMPR73[6] , \R_DATA_TEMPR73[5] , \R_DATA_TEMPR73[4] , 
        \R_DATA_TEMPR73[3] , \R_DATA_TEMPR73[2] , \R_DATA_TEMPR73[1] , 
        \R_DATA_TEMPR73[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[73][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[18] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[18] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1340 (.A(OR4_1494_Y), .B(OR4_107_Y), .C(OR4_309_Y), .D(
        OR4_1578_Y), .Y(OR4_1340_Y));
    OR4 OR4_656 (.A(OR4_411_Y), .B(OR4_1157_Y), .C(OR4_73_Y), .D(
        OR4_1093_Y), .Y(OR4_656_Y));
    OR4 OR4_1117 (.A(\R_DATA_TEMPR16[8] ), .B(\R_DATA_TEMPR17[8] ), .C(
        \R_DATA_TEMPR18[8] ), .D(\R_DATA_TEMPR19[8] ), .Y(OR4_1117_Y));
    OR4 OR4_440 (.A(OR4_1441_Y), .B(OR4_906_Y), .C(OR4_1461_Y), .D(
        OR4_841_Y), .Y(OR4_440_Y));
    OR4 OR4_1266 (.A(OR4_1321_Y), .B(OR4_1042_Y), .C(OR4_764_Y), .D(
        OR4_1277_Y), .Y(OR4_1266_Y));
    OR4 OR4_293 (.A(\R_DATA_TEMPR28[1] ), .B(\R_DATA_TEMPR29[1] ), .C(
        \R_DATA_TEMPR30[1] ), .D(\R_DATA_TEMPR31[1] ), .Y(OR4_293_Y));
    OR4 OR4_388 (.A(OR4_229_Y), .B(OR4_757_Y), .C(OR4_400_Y), .D(
        OR4_396_Y), .Y(OR4_388_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%83%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R83C0 (.A_DOUT({
        \R_DATA_TEMPR83[39] , \R_DATA_TEMPR83[38] , 
        \R_DATA_TEMPR83[37] , \R_DATA_TEMPR83[36] , 
        \R_DATA_TEMPR83[35] , \R_DATA_TEMPR83[34] , 
        \R_DATA_TEMPR83[33] , \R_DATA_TEMPR83[32] , 
        \R_DATA_TEMPR83[31] , \R_DATA_TEMPR83[30] , 
        \R_DATA_TEMPR83[29] , \R_DATA_TEMPR83[28] , 
        \R_DATA_TEMPR83[27] , \R_DATA_TEMPR83[26] , 
        \R_DATA_TEMPR83[25] , \R_DATA_TEMPR83[24] , 
        \R_DATA_TEMPR83[23] , \R_DATA_TEMPR83[22] , 
        \R_DATA_TEMPR83[21] , \R_DATA_TEMPR83[20] }), .B_DOUT({
        \R_DATA_TEMPR83[19] , \R_DATA_TEMPR83[18] , 
        \R_DATA_TEMPR83[17] , \R_DATA_TEMPR83[16] , 
        \R_DATA_TEMPR83[15] , \R_DATA_TEMPR83[14] , 
        \R_DATA_TEMPR83[13] , \R_DATA_TEMPR83[12] , 
        \R_DATA_TEMPR83[11] , \R_DATA_TEMPR83[10] , 
        \R_DATA_TEMPR83[9] , \R_DATA_TEMPR83[8] , \R_DATA_TEMPR83[7] , 
        \R_DATA_TEMPR83[6] , \R_DATA_TEMPR83[5] , \R_DATA_TEMPR83[4] , 
        \R_DATA_TEMPR83[3] , \R_DATA_TEMPR83[2] , \R_DATA_TEMPR83[1] , 
        \R_DATA_TEMPR83[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[83][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[20] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[20] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_115 (.A(OR4_667_Y), .B(OR4_1189_Y), .C(OR4_694_Y), .D(
        OR4_205_Y), .Y(OR4_115_Y));
    OR4 OR4_66 (.A(OR4_522_Y), .B(OR4_363_Y), .C(OR4_481_Y), .D(
        OR4_94_Y), .Y(OR4_66_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%56%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R56C0 (.A_DOUT({
        \R_DATA_TEMPR56[39] , \R_DATA_TEMPR56[38] , 
        \R_DATA_TEMPR56[37] , \R_DATA_TEMPR56[36] , 
        \R_DATA_TEMPR56[35] , \R_DATA_TEMPR56[34] , 
        \R_DATA_TEMPR56[33] , \R_DATA_TEMPR56[32] , 
        \R_DATA_TEMPR56[31] , \R_DATA_TEMPR56[30] , 
        \R_DATA_TEMPR56[29] , \R_DATA_TEMPR56[28] , 
        \R_DATA_TEMPR56[27] , \R_DATA_TEMPR56[26] , 
        \R_DATA_TEMPR56[25] , \R_DATA_TEMPR56[24] , 
        \R_DATA_TEMPR56[23] , \R_DATA_TEMPR56[22] , 
        \R_DATA_TEMPR56[21] , \R_DATA_TEMPR56[20] }), .B_DOUT({
        \R_DATA_TEMPR56[19] , \R_DATA_TEMPR56[18] , 
        \R_DATA_TEMPR56[17] , \R_DATA_TEMPR56[16] , 
        \R_DATA_TEMPR56[15] , \R_DATA_TEMPR56[14] , 
        \R_DATA_TEMPR56[13] , \R_DATA_TEMPR56[12] , 
        \R_DATA_TEMPR56[11] , \R_DATA_TEMPR56[10] , 
        \R_DATA_TEMPR56[9] , \R_DATA_TEMPR56[8] , \R_DATA_TEMPR56[7] , 
        \R_DATA_TEMPR56[6] , \R_DATA_TEMPR56[5] , \R_DATA_TEMPR56[4] , 
        \R_DATA_TEMPR56[3] , \R_DATA_TEMPR56[2] , \R_DATA_TEMPR56[1] , 
        \R_DATA_TEMPR56[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[56][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[14] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[14] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1368 (.A(\R_DATA_TEMPR44[32] ), .B(\R_DATA_TEMPR45[32] ), 
        .C(\R_DATA_TEMPR46[32] ), .D(\R_DATA_TEMPR47[32] ), .Y(
        OR4_1368_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[24]  (.A(CFG3_13_Y), .B(
        CFG3_7_Y), .Y(\BLKX2[24] ));
    OR4 OR4_998 (.A(\R_DATA_TEMPR0[24] ), .B(\R_DATA_TEMPR1[24] ), .C(
        \R_DATA_TEMPR2[24] ), .D(\R_DATA_TEMPR3[24] ), .Y(OR4_998_Y));
    OR4 OR4_417 (.A(\R_DATA_TEMPR12[38] ), .B(\R_DATA_TEMPR13[38] ), 
        .C(\R_DATA_TEMPR14[38] ), .D(\R_DATA_TEMPR15[38] ), .Y(
        OR4_417_Y));
    OR4 OR4_433 (.A(\R_DATA_TEMPR104[10] ), .B(\R_DATA_TEMPR105[10] ), 
        .C(\R_DATA_TEMPR106[10] ), .D(\R_DATA_TEMPR107[10] ), .Y(
        OR4_433_Y));
    OR4 OR4_631 (.A(\R_DATA_TEMPR52[14] ), .B(\R_DATA_TEMPR53[14] ), 
        .C(\R_DATA_TEMPR54[14] ), .D(\R_DATA_TEMPR55[14] ), .Y(
        OR4_631_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%46%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R46C0 (.A_DOUT({
        \R_DATA_TEMPR46[39] , \R_DATA_TEMPR46[38] , 
        \R_DATA_TEMPR46[37] , \R_DATA_TEMPR46[36] , 
        \R_DATA_TEMPR46[35] , \R_DATA_TEMPR46[34] , 
        \R_DATA_TEMPR46[33] , \R_DATA_TEMPR46[32] , 
        \R_DATA_TEMPR46[31] , \R_DATA_TEMPR46[30] , 
        \R_DATA_TEMPR46[29] , \R_DATA_TEMPR46[28] , 
        \R_DATA_TEMPR46[27] , \R_DATA_TEMPR46[26] , 
        \R_DATA_TEMPR46[25] , \R_DATA_TEMPR46[24] , 
        \R_DATA_TEMPR46[23] , \R_DATA_TEMPR46[22] , 
        \R_DATA_TEMPR46[21] , \R_DATA_TEMPR46[20] }), .B_DOUT({
        \R_DATA_TEMPR46[19] , \R_DATA_TEMPR46[18] , 
        \R_DATA_TEMPR46[17] , \R_DATA_TEMPR46[16] , 
        \R_DATA_TEMPR46[15] , \R_DATA_TEMPR46[14] , 
        \R_DATA_TEMPR46[13] , \R_DATA_TEMPR46[12] , 
        \R_DATA_TEMPR46[11] , \R_DATA_TEMPR46[10] , 
        \R_DATA_TEMPR46[9] , \R_DATA_TEMPR46[8] , \R_DATA_TEMPR46[7] , 
        \R_DATA_TEMPR46[6] , \R_DATA_TEMPR46[5] , \R_DATA_TEMPR46[4] , 
        \R_DATA_TEMPR46[3] , \R_DATA_TEMPR46[2] , \R_DATA_TEMPR46[1] , 
        \R_DATA_TEMPR46[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[46][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[11] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[11] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_365 (.A(OR4_1311_Y), .B(OR4_1614_Y), .C(OR4_1054_Y), .D(
        OR4_289_Y), .Y(OR4_365_Y));
    OR4 OR4_238 (.A(\R_DATA_TEMPR4[3] ), .B(\R_DATA_TEMPR5[3] ), .C(
        \R_DATA_TEMPR6[3] ), .D(\R_DATA_TEMPR7[3] ), .Y(OR4_238_Y));
    OR2 OR2_8 (.A(\R_DATA_TEMPR84[1] ), .B(\R_DATA_TEMPR85[1] ), .Y(
        OR2_8_Y));
    OR4 OR4_189 (.A(\R_DATA_TEMPR100[10] ), .B(\R_DATA_TEMPR101[10] ), 
        .C(\R_DATA_TEMPR102[10] ), .D(\R_DATA_TEMPR103[10] ), .Y(
        OR4_189_Y));
    OR4 OR4_0 (.A(\R_DATA_TEMPR80[11] ), .B(\R_DATA_TEMPR81[11] ), .C(
        \R_DATA_TEMPR82[11] ), .D(\R_DATA_TEMPR83[11] ), .Y(OR4_0_Y));
    OR4 OR4_1473 (.A(\R_DATA_TEMPR8[29] ), .B(\R_DATA_TEMPR9[29] ), .C(
        \R_DATA_TEMPR10[29] ), .D(\R_DATA_TEMPR11[29] ), .Y(OR4_1473_Y)
        );
    OR4 OR4_207 (.A(\R_DATA_TEMPR120[39] ), .B(\R_DATA_TEMPR121[39] ), 
        .C(\R_DATA_TEMPR122[39] ), .D(\R_DATA_TEMPR123[39] ), .Y(
        OR4_207_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%68%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R68C0 (.A_DOUT({
        \R_DATA_TEMPR68[39] , \R_DATA_TEMPR68[38] , 
        \R_DATA_TEMPR68[37] , \R_DATA_TEMPR68[36] , 
        \R_DATA_TEMPR68[35] , \R_DATA_TEMPR68[34] , 
        \R_DATA_TEMPR68[33] , \R_DATA_TEMPR68[32] , 
        \R_DATA_TEMPR68[31] , \R_DATA_TEMPR68[30] , 
        \R_DATA_TEMPR68[29] , \R_DATA_TEMPR68[28] , 
        \R_DATA_TEMPR68[27] , \R_DATA_TEMPR68[26] , 
        \R_DATA_TEMPR68[25] , \R_DATA_TEMPR68[24] , 
        \R_DATA_TEMPR68[23] , \R_DATA_TEMPR68[22] , 
        \R_DATA_TEMPR68[21] , \R_DATA_TEMPR68[20] }), .B_DOUT({
        \R_DATA_TEMPR68[19] , \R_DATA_TEMPR68[18] , 
        \R_DATA_TEMPR68[17] , \R_DATA_TEMPR68[16] , 
        \R_DATA_TEMPR68[15] , \R_DATA_TEMPR68[14] , 
        \R_DATA_TEMPR68[13] , \R_DATA_TEMPR68[12] , 
        \R_DATA_TEMPR68[11] , \R_DATA_TEMPR68[10] , 
        \R_DATA_TEMPR68[9] , \R_DATA_TEMPR68[8] , \R_DATA_TEMPR68[7] , 
        \R_DATA_TEMPR68[6] , \R_DATA_TEMPR68[5] , \R_DATA_TEMPR68[4] , 
        \R_DATA_TEMPR68[3] , \R_DATA_TEMPR68[2] , \R_DATA_TEMPR68[1] , 
        \R_DATA_TEMPR68[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[68][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[17] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[17] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_215 (.A(OR4_358_Y), .B(OR4_1248_Y), .C(OR4_247_Y), .D(
        OR4_1012_Y), .Y(OR4_215_Y));
    OR4 OR4_1245 (.A(\R_DATA_TEMPR120[23] ), .B(\R_DATA_TEMPR121[23] ), 
        .C(\R_DATA_TEMPR122[23] ), .D(\R_DATA_TEMPR123[23] ), .Y(
        OR4_1245_Y));
    OR4 OR4_107 (.A(\R_DATA_TEMPR116[0] ), .B(\R_DATA_TEMPR117[0] ), 
        .C(\R_DATA_TEMPR118[0] ), .D(\R_DATA_TEMPR119[0] ), .Y(
        OR4_107_Y));
    OR4 OR4_1002 (.A(OR4_1075_Y), .B(OR4_858_Y), .C(OR4_1403_Y), .D(
        OR4_212_Y), .Y(OR4_1002_Y));
    OR4 OR4_1069 (.A(OR4_1605_Y), .B(OR4_225_Y), .C(OR4_1371_Y), .D(
        OR4_1095_Y), .Y(OR4_1069_Y));
    OR4 OR4_1595 (.A(\R_DATA_TEMPR32[8] ), .B(\R_DATA_TEMPR33[8] ), .C(
        \R_DATA_TEMPR34[8] ), .D(\R_DATA_TEMPR35[8] ), .Y(OR4_1595_Y));
    OR4 OR4_812 (.A(\R_DATA_TEMPR32[37] ), .B(\R_DATA_TEMPR33[37] ), 
        .C(\R_DATA_TEMPR34[37] ), .D(\R_DATA_TEMPR35[37] ), .Y(
        OR4_812_Y));
    OR4 OR4_277 (.A(\R_DATA_TEMPR0[37] ), .B(\R_DATA_TEMPR1[37] ), .C(
        \R_DATA_TEMPR2[37] ), .D(\R_DATA_TEMPR3[37] ), .Y(OR4_277_Y));
    OR4 OR4_1541 (.A(\R_DATA_TEMPR4[9] ), .B(\R_DATA_TEMPR5[9] ), .C(
        \R_DATA_TEMPR6[9] ), .D(\R_DATA_TEMPR7[9] ), .Y(OR4_1541_Y));
    OR4 OR4_698 (.A(\R_DATA_TEMPR32[13] ), .B(\R_DATA_TEMPR33[13] ), 
        .C(\R_DATA_TEMPR34[13] ), .D(\R_DATA_TEMPR35[13] ), .Y(
        OR4_698_Y));
    OR4 OR4_95 (.A(\R_DATA_TEMPR112[18] ), .B(\R_DATA_TEMPR113[18] ), 
        .C(\R_DATA_TEMPR114[18] ), .D(\R_DATA_TEMPR115[18] ), .Y(
        OR4_95_Y));
    OR4 OR4_1538 (.A(\R_DATA_TEMPR56[10] ), .B(\R_DATA_TEMPR57[10] ), 
        .C(\R_DATA_TEMPR58[10] ), .D(\R_DATA_TEMPR59[10] ), .Y(
        OR4_1538_Y));
    OR2 OR2_22 (.A(\R_DATA_TEMPR84[11] ), .B(\R_DATA_TEMPR85[11] ), .Y(
        OR2_22_Y));
    OR4 OR4_177 (.A(\R_DATA_TEMPR92[26] ), .B(\R_DATA_TEMPR93[26] ), 
        .C(\R_DATA_TEMPR94[26] ), .D(\R_DATA_TEMPR95[26] ), .Y(
        OR4_177_Y));
    OR4 \OR4_R_DATA[34]  (.A(OR4_310_Y), .B(OR4_1362_Y), .C(OR4_531_Y), 
        .D(OR4_1229_Y), .Y(R_DATA[34]));
    OR4 OR4_981 (.A(\R_DATA_TEMPR76[30] ), .B(\R_DATA_TEMPR77[30] ), 
        .C(\R_DATA_TEMPR78[30] ), .D(\R_DATA_TEMPR79[30] ), .Y(
        OR4_981_Y));
    OR4 OR4_1296 (.A(\R_DATA_TEMPR116[26] ), .B(\R_DATA_TEMPR117[26] ), 
        .C(\R_DATA_TEMPR118[26] ), .D(\R_DATA_TEMPR119[26] ), .Y(
        OR4_1296_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[14]  (.A(CFG3_1_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[14] ));
    OR4 OR4_762 (.A(\R_DATA_TEMPR80[25] ), .B(\R_DATA_TEMPR81[25] ), 
        .C(\R_DATA_TEMPR82[25] ), .D(\R_DATA_TEMPR83[25] ), .Y(
        OR4_762_Y));
    OR4 OR4_349 (.A(\R_DATA_TEMPR24[19] ), .B(\R_DATA_TEMPR25[19] ), 
        .C(\R_DATA_TEMPR26[19] ), .D(\R_DATA_TEMPR27[19] ), .Y(
        OR4_349_Y));
    OR4 OR4_1239 (.A(\R_DATA_TEMPR100[23] ), .B(\R_DATA_TEMPR101[23] ), 
        .C(\R_DATA_TEMPR102[23] ), .D(\R_DATA_TEMPR103[23] ), .Y(
        OR4_1239_Y));
    OR4 OR4_692 (.A(\R_DATA_TEMPR20[19] ), .B(\R_DATA_TEMPR21[19] ), 
        .C(\R_DATA_TEMPR22[19] ), .D(\R_DATA_TEMPR23[19] ), .Y(
        OR4_692_Y));
    OR4 OR4_1210 (.A(\R_DATA_TEMPR64[1] ), .B(\R_DATA_TEMPR65[1] ), .C(
        \R_DATA_TEMPR66[1] ), .D(\R_DATA_TEMPR67[1] ), .Y(OR4_1210_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[31]  (.A(CFG3_21_Y), .B(
        CFG3_3_Y), .Y(\BLKY2[31] ));
    OR4 OR4_703 (.A(\R_DATA_TEMPR64[27] ), .B(\R_DATA_TEMPR65[27] ), 
        .C(\R_DATA_TEMPR66[27] ), .D(\R_DATA_TEMPR67[27] ), .Y(
        OR4_703_Y));
    OR4 OR4_223 (.A(OR4_285_Y), .B(OR4_1601_Y), .C(OR4_391_Y), .D(
        OR4_213_Y), .Y(OR4_223_Y));
    OR4 OR4_1398 (.A(\R_DATA_TEMPR48[0] ), .B(\R_DATA_TEMPR49[0] ), .C(
        \R_DATA_TEMPR50[0] ), .D(\R_DATA_TEMPR51[0] ), .Y(OR4_1398_Y));
    OR4 OR4_966 (.A(\R_DATA_TEMPR76[32] ), .B(\R_DATA_TEMPR77[32] ), 
        .C(\R_DATA_TEMPR78[32] ), .D(\R_DATA_TEMPR79[32] ), .Y(
        OR4_966_Y));
    OR4 OR4_204 (.A(\R_DATA_TEMPR80[9] ), .B(\R_DATA_TEMPR81[9] ), .C(
        \R_DATA_TEMPR82[9] ), .D(\R_DATA_TEMPR83[9] ), .Y(OR4_204_Y));
    OR4 OR4_354 (.A(OR4_1394_Y), .B(OR4_1113_Y), .C(OR4_833_Y), .D(
        OR4_316_Y), .Y(OR4_354_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%29%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C0 (.A_DOUT({
        \R_DATA_TEMPR29[39] , \R_DATA_TEMPR29[38] , 
        \R_DATA_TEMPR29[37] , \R_DATA_TEMPR29[36] , 
        \R_DATA_TEMPR29[35] , \R_DATA_TEMPR29[34] , 
        \R_DATA_TEMPR29[33] , \R_DATA_TEMPR29[32] , 
        \R_DATA_TEMPR29[31] , \R_DATA_TEMPR29[30] , 
        \R_DATA_TEMPR29[29] , \R_DATA_TEMPR29[28] , 
        \R_DATA_TEMPR29[27] , \R_DATA_TEMPR29[26] , 
        \R_DATA_TEMPR29[25] , \R_DATA_TEMPR29[24] , 
        \R_DATA_TEMPR29[23] , \R_DATA_TEMPR29[22] , 
        \R_DATA_TEMPR29[21] , \R_DATA_TEMPR29[20] }), .B_DOUT({
        \R_DATA_TEMPR29[19] , \R_DATA_TEMPR29[18] , 
        \R_DATA_TEMPR29[17] , \R_DATA_TEMPR29[16] , 
        \R_DATA_TEMPR29[15] , \R_DATA_TEMPR29[14] , 
        \R_DATA_TEMPR29[13] , \R_DATA_TEMPR29[12] , 
        \R_DATA_TEMPR29[11] , \R_DATA_TEMPR29[10] , 
        \R_DATA_TEMPR29[9] , \R_DATA_TEMPR29[8] , \R_DATA_TEMPR29[7] , 
        \R_DATA_TEMPR29[6] , \R_DATA_TEMPR29[5] , \R_DATA_TEMPR29[4] , 
        \R_DATA_TEMPR29[3] , \R_DATA_TEMPR29[2] , \R_DATA_TEMPR29[1] , 
        \R_DATA_TEMPR29[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR2 OR2_19 (.A(\R_DATA_TEMPR84[9] ), .B(\R_DATA_TEMPR85[9] ), .Y(
        OR2_19_Y));
    OR4 OR4_1517 (.A(\R_DATA_TEMPR20[14] ), .B(\R_DATA_TEMPR21[14] ), 
        .C(\R_DATA_TEMPR22[14] ), .D(\R_DATA_TEMPR23[14] ), .Y(
        OR4_1517_Y));
    OR4 OR4_773 (.A(OR4_438_Y), .B(OR4_1570_Y), .C(OR4_1625_Y), .D(
        OR4_1175_Y), .Y(OR4_773_Y));
    OR4 OR4_665 (.A(OR4_856_Y), .B(OR4_1108_Y), .C(OR4_1305_Y), .D(
        OR4_879_Y), .Y(OR4_665_Y));
    OR4 OR4_413 (.A(\R_DATA_TEMPR56[36] ), .B(\R_DATA_TEMPR57[36] ), 
        .C(\R_DATA_TEMPR58[36] ), .D(\R_DATA_TEMPR59[36] ), .Y(
        OR4_413_Y));
    OR4 OR4_611 (.A(\R_DATA_TEMPR116[9] ), .B(\R_DATA_TEMPR117[9] ), 
        .C(\R_DATA_TEMPR118[9] ), .D(\R_DATA_TEMPR119[9] ), .Y(
        OR4_611_Y));
    OR4 OR4_1312 (.A(\R_DATA_TEMPR96[21] ), .B(\R_DATA_TEMPR97[21] ), 
        .C(\R_DATA_TEMPR98[21] ), .D(\R_DATA_TEMPR99[21] ), .Y(
        OR4_1312_Y));
    OR4 OR4_1082 (.A(\R_DATA_TEMPR44[6] ), .B(\R_DATA_TEMPR45[6] ), .C(
        \R_DATA_TEMPR46[6] ), .D(\R_DATA_TEMPR47[6] ), .Y(OR4_1082_Y));
    OR4 OR4_928 (.A(\R_DATA_TEMPR104[8] ), .B(\R_DATA_TEMPR105[8] ), 
        .C(\R_DATA_TEMPR106[8] ), .D(\R_DATA_TEMPR107[8] ), .Y(
        OR4_928_Y));
    OR4 OR4_151 (.A(OR4_1228_Y), .B(OR2_25_Y), .C(\R_DATA_TEMPR86[33] )
        , .D(\R_DATA_TEMPR87[33] ), .Y(OR4_151_Y));
    OR4 OR4_274 (.A(\R_DATA_TEMPR120[1] ), .B(\R_DATA_TEMPR121[1] ), 
        .C(\R_DATA_TEMPR122[1] ), .D(\R_DATA_TEMPR123[1] ), .Y(
        OR4_274_Y));
    OR4 OR4_218 (.A(\R_DATA_TEMPR64[19] ), .B(\R_DATA_TEMPR65[19] ), 
        .C(\R_DATA_TEMPR66[19] ), .D(\R_DATA_TEMPR67[19] ), .Y(
        OR4_218_Y));
    OR4 OR4_1554 (.A(OR4_1053_Y), .B(OR4_715_Y), .C(OR4_451_Y), .D(
        OR4_533_Y), .Y(OR4_1554_Y));
    OR4 OR4_1212 (.A(\R_DATA_TEMPR4[29] ), .B(\R_DATA_TEMPR5[29] ), .C(
        \R_DATA_TEMPR6[29] ), .D(\R_DATA_TEMPR7[29] ), .Y(OR4_1212_Y));
    OR4 \OR4_R_DATA[22]  (.A(OR4_1038_Y), .B(OR4_991_Y), .C(OR4_772_Y), 
        .D(OR4_38_Y), .Y(R_DATA[22]));
    OR4 OR4_60 (.A(\R_DATA_TEMPR60[3] ), .B(\R_DATA_TEMPR61[3] ), .C(
        \R_DATA_TEMPR62[3] ), .D(\R_DATA_TEMPR63[3] ), .Y(OR4_60_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%111%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R111C0 (.A_DOUT({
        \R_DATA_TEMPR111[39] , \R_DATA_TEMPR111[38] , 
        \R_DATA_TEMPR111[37] , \R_DATA_TEMPR111[36] , 
        \R_DATA_TEMPR111[35] , \R_DATA_TEMPR111[34] , 
        \R_DATA_TEMPR111[33] , \R_DATA_TEMPR111[32] , 
        \R_DATA_TEMPR111[31] , \R_DATA_TEMPR111[30] , 
        \R_DATA_TEMPR111[29] , \R_DATA_TEMPR111[28] , 
        \R_DATA_TEMPR111[27] , \R_DATA_TEMPR111[26] , 
        \R_DATA_TEMPR111[25] , \R_DATA_TEMPR111[24] , 
        \R_DATA_TEMPR111[23] , \R_DATA_TEMPR111[22] , 
        \R_DATA_TEMPR111[21] , \R_DATA_TEMPR111[20] }), .B_DOUT({
        \R_DATA_TEMPR111[19] , \R_DATA_TEMPR111[18] , 
        \R_DATA_TEMPR111[17] , \R_DATA_TEMPR111[16] , 
        \R_DATA_TEMPR111[15] , \R_DATA_TEMPR111[14] , 
        \R_DATA_TEMPR111[13] , \R_DATA_TEMPR111[12] , 
        \R_DATA_TEMPR111[11] , \R_DATA_TEMPR111[10] , 
        \R_DATA_TEMPR111[9] , \R_DATA_TEMPR111[8] , 
        \R_DATA_TEMPR111[7] , \R_DATA_TEMPR111[6] , 
        \R_DATA_TEMPR111[5] , \R_DATA_TEMPR111[4] , 
        \R_DATA_TEMPR111[3] , \R_DATA_TEMPR111[2] , 
        \R_DATA_TEMPR111[1] , \R_DATA_TEMPR111[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[111][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[27] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[27] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1355 (.A(\R_DATA_TEMPR112[12] ), .B(\R_DATA_TEMPR113[12] ), 
        .C(\R_DATA_TEMPR114[12] ), .D(\R_DATA_TEMPR115[12] ), .Y(
        OR4_1355_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%98%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R98C0 (.A_DOUT({
        \R_DATA_TEMPR98[39] , \R_DATA_TEMPR98[38] , 
        \R_DATA_TEMPR98[37] , \R_DATA_TEMPR98[36] , 
        \R_DATA_TEMPR98[35] , \R_DATA_TEMPR98[34] , 
        \R_DATA_TEMPR98[33] , \R_DATA_TEMPR98[32] , 
        \R_DATA_TEMPR98[31] , \R_DATA_TEMPR98[30] , 
        \R_DATA_TEMPR98[29] , \R_DATA_TEMPR98[28] , 
        \R_DATA_TEMPR98[27] , \R_DATA_TEMPR98[26] , 
        \R_DATA_TEMPR98[25] , \R_DATA_TEMPR98[24] , 
        \R_DATA_TEMPR98[23] , \R_DATA_TEMPR98[22] , 
        \R_DATA_TEMPR98[21] , \R_DATA_TEMPR98[20] }), .B_DOUT({
        \R_DATA_TEMPR98[19] , \R_DATA_TEMPR98[18] , 
        \R_DATA_TEMPR98[17] , \R_DATA_TEMPR98[16] , 
        \R_DATA_TEMPR98[15] , \R_DATA_TEMPR98[14] , 
        \R_DATA_TEMPR98[13] , \R_DATA_TEMPR98[12] , 
        \R_DATA_TEMPR98[11] , \R_DATA_TEMPR98[10] , 
        \R_DATA_TEMPR98[9] , \R_DATA_TEMPR98[8] , \R_DATA_TEMPR98[7] , 
        \R_DATA_TEMPR98[6] , \R_DATA_TEMPR98[5] , \R_DATA_TEMPR98[4] , 
        \R_DATA_TEMPR98[3] , \R_DATA_TEMPR98[2] , \R_DATA_TEMPR98[1] , 
        \R_DATA_TEMPR98[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[98][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[24] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[24] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_531 (.A(OR4_797_Y), .B(OR4_624_Y), .C(OR4_16_Y), .D(
        OR4_550_Y), .Y(OR4_531_Y));
    OR4 OR4_1414 (.A(\R_DATA_TEMPR28[8] ), .B(\R_DATA_TEMPR29[8] ), .C(
        \R_DATA_TEMPR30[8] ), .D(\R_DATA_TEMPR31[8] ), .Y(OR4_1414_Y));
    OR4 OR4_1099 (.A(\R_DATA_TEMPR36[13] ), .B(\R_DATA_TEMPR37[13] ), 
        .C(\R_DATA_TEMPR38[13] ), .D(\R_DATA_TEMPR39[13] ), .Y(
        OR4_1099_Y));
    OR4 OR4_895 (.A(\R_DATA_TEMPR20[5] ), .B(\R_DATA_TEMPR21[5] ), .C(
        \R_DATA_TEMPR22[5] ), .D(\R_DATA_TEMPR23[5] ), .Y(OR4_895_Y));
    OR4 OR4_67 (.A(\R_DATA_TEMPR48[30] ), .B(\R_DATA_TEMPR49[30] ), .C(
        \R_DATA_TEMPR50[30] ), .D(\R_DATA_TEMPR51[30] ), .Y(OR4_67_Y));
    OR4 OR4_785 (.A(\R_DATA_TEMPR20[22] ), .B(\R_DATA_TEMPR21[22] ), 
        .C(\R_DATA_TEMPR22[22] ), .D(\R_DATA_TEMPR23[22] ), .Y(
        OR4_785_Y));
    OR4 OR4_687 (.A(\R_DATA_TEMPR28[29] ), .B(\R_DATA_TEMPR29[29] ), 
        .C(\R_DATA_TEMPR30[29] ), .D(\R_DATA_TEMPR31[29] ), .Y(
        OR4_687_Y));
    OR4 OR4_305 (.A(\R_DATA_TEMPR124[37] ), .B(\R_DATA_TEMPR125[37] ), 
        .C(\R_DATA_TEMPR126[37] ), .D(\R_DATA_TEMPR127[37] ), .Y(
        OR4_305_Y));
    OR4 OR4_451 (.A(OR4_1483_Y), .B(OR4_1170_Y), .C(OR4_1141_Y), .D(
        OR4_320_Y), .Y(OR4_451_Y));
    OR4 OR4_1214 (.A(\R_DATA_TEMPR52[33] ), .B(\R_DATA_TEMPR53[33] ), 
        .C(\R_DATA_TEMPR54[33] ), .D(\R_DATA_TEMPR55[33] ), .Y(
        OR4_1214_Y));
    OR4 OR4_786 (.A(\R_DATA_TEMPR0[36] ), .B(\R_DATA_TEMPR1[36] ), .C(
        \R_DATA_TEMPR2[36] ), .D(\R_DATA_TEMPR3[36] ), .Y(OR4_786_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%105%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R105C0 (.A_DOUT({
        \R_DATA_TEMPR105[39] , \R_DATA_TEMPR105[38] , 
        \R_DATA_TEMPR105[37] , \R_DATA_TEMPR105[36] , 
        \R_DATA_TEMPR105[35] , \R_DATA_TEMPR105[34] , 
        \R_DATA_TEMPR105[33] , \R_DATA_TEMPR105[32] , 
        \R_DATA_TEMPR105[31] , \R_DATA_TEMPR105[30] , 
        \R_DATA_TEMPR105[29] , \R_DATA_TEMPR105[28] , 
        \R_DATA_TEMPR105[27] , \R_DATA_TEMPR105[26] , 
        \R_DATA_TEMPR105[25] , \R_DATA_TEMPR105[24] , 
        \R_DATA_TEMPR105[23] , \R_DATA_TEMPR105[22] , 
        \R_DATA_TEMPR105[21] , \R_DATA_TEMPR105[20] }), .B_DOUT({
        \R_DATA_TEMPR105[19] , \R_DATA_TEMPR105[18] , 
        \R_DATA_TEMPR105[17] , \R_DATA_TEMPR105[16] , 
        \R_DATA_TEMPR105[15] , \R_DATA_TEMPR105[14] , 
        \R_DATA_TEMPR105[13] , \R_DATA_TEMPR105[12] , 
        \R_DATA_TEMPR105[11] , \R_DATA_TEMPR105[10] , 
        \R_DATA_TEMPR105[9] , \R_DATA_TEMPR105[8] , 
        \R_DATA_TEMPR105[7] , \R_DATA_TEMPR105[6] , 
        \R_DATA_TEMPR105[5] , \R_DATA_TEMPR105[4] , 
        \R_DATA_TEMPR105[3] , \R_DATA_TEMPR105[2] , 
        \R_DATA_TEMPR105[1] , \R_DATA_TEMPR105[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[105][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[26] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[26] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1528 (.A(\R_DATA_TEMPR116[23] ), .B(\R_DATA_TEMPR117[23] ), 
        .C(\R_DATA_TEMPR118[23] ), .D(\R_DATA_TEMPR119[23] ), .Y(
        OR4_1528_Y));
    OR4 OR4_1503 (.A(OR4_377_Y), .B(OR4_632_Y), .C(OR4_129_Y), .D(
        OR4_1515_Y), .Y(OR4_1503_Y));
    OR4 OR4_458 (.A(\R_DATA_TEMPR48[35] ), .B(\R_DATA_TEMPR49[35] ), 
        .C(\R_DATA_TEMPR50[35] ), .D(\R_DATA_TEMPR51[35] ), .Y(
        OR4_458_Y));
    OR4 OR4_1173 (.A(\R_DATA_TEMPR116[12] ), .B(\R_DATA_TEMPR117[12] ), 
        .C(\R_DATA_TEMPR118[12] ), .D(\R_DATA_TEMPR119[12] ), .Y(
        OR4_1173_Y));
    OR4 OR4_628 (.A(\R_DATA_TEMPR40[6] ), .B(\R_DATA_TEMPR41[6] ), .C(
        \R_DATA_TEMPR42[6] ), .D(\R_DATA_TEMPR43[6] ), .Y(OR4_628_Y));
    OR4 OR4_375 (.A(OR4_661_Y), .B(OR4_1239_Y), .C(OR4_401_Y), .D(
        OR4_651_Y), .Y(OR4_375_Y));
    OR4 OR4_1317 (.A(\R_DATA_TEMPR56[35] ), .B(\R_DATA_TEMPR57[35] ), 
        .C(\R_DATA_TEMPR58[35] ), .D(\R_DATA_TEMPR59[35] ), .Y(
        OR4_1317_Y));
    OR4 OR4_749 (.A(\R_DATA_TEMPR80[10] ), .B(\R_DATA_TEMPR81[10] ), 
        .C(\R_DATA_TEMPR82[10] ), .D(\R_DATA_TEMPR83[10] ), .Y(
        OR4_749_Y));
    OR4 OR4_1229 (.A(OR4_46_Y), .B(OR4_1172_Y), .C(OR4_1232_Y), .D(
        OR4_134_Y), .Y(OR4_1229_Y));
    OR4 OR4_660 (.A(\R_DATA_TEMPR108[1] ), .B(\R_DATA_TEMPR109[1] ), 
        .C(\R_DATA_TEMPR110[1] ), .D(\R_DATA_TEMPR111[1] ), .Y(
        OR4_660_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%25%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C0 (.A_DOUT({
        \R_DATA_TEMPR25[39] , \R_DATA_TEMPR25[38] , 
        \R_DATA_TEMPR25[37] , \R_DATA_TEMPR25[36] , 
        \R_DATA_TEMPR25[35] , \R_DATA_TEMPR25[34] , 
        \R_DATA_TEMPR25[33] , \R_DATA_TEMPR25[32] , 
        \R_DATA_TEMPR25[31] , \R_DATA_TEMPR25[30] , 
        \R_DATA_TEMPR25[29] , \R_DATA_TEMPR25[28] , 
        \R_DATA_TEMPR25[27] , \R_DATA_TEMPR25[26] , 
        \R_DATA_TEMPR25[25] , \R_DATA_TEMPR25[24] , 
        \R_DATA_TEMPR25[23] , \R_DATA_TEMPR25[22] , 
        \R_DATA_TEMPR25[21] , \R_DATA_TEMPR25[20] }), .B_DOUT({
        \R_DATA_TEMPR25[19] , \R_DATA_TEMPR25[18] , 
        \R_DATA_TEMPR25[17] , \R_DATA_TEMPR25[16] , 
        \R_DATA_TEMPR25[15] , \R_DATA_TEMPR25[14] , 
        \R_DATA_TEMPR25[13] , \R_DATA_TEMPR25[12] , 
        \R_DATA_TEMPR25[11] , \R_DATA_TEMPR25[10] , 
        \R_DATA_TEMPR25[9] , \R_DATA_TEMPR25[8] , \R_DATA_TEMPR25[7] , 
        \R_DATA_TEMPR25[6] , \R_DATA_TEMPR25[5] , \R_DATA_TEMPR25[4] , 
        \R_DATA_TEMPR25[3] , \R_DATA_TEMPR25[2] , \R_DATA_TEMPR25[1] , 
        \R_DATA_TEMPR25[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%67%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R67C0 (.A_DOUT({
        \R_DATA_TEMPR67[39] , \R_DATA_TEMPR67[38] , 
        \R_DATA_TEMPR67[37] , \R_DATA_TEMPR67[36] , 
        \R_DATA_TEMPR67[35] , \R_DATA_TEMPR67[34] , 
        \R_DATA_TEMPR67[33] , \R_DATA_TEMPR67[32] , 
        \R_DATA_TEMPR67[31] , \R_DATA_TEMPR67[30] , 
        \R_DATA_TEMPR67[29] , \R_DATA_TEMPR67[28] , 
        \R_DATA_TEMPR67[27] , \R_DATA_TEMPR67[26] , 
        \R_DATA_TEMPR67[25] , \R_DATA_TEMPR67[24] , 
        \R_DATA_TEMPR67[23] , \R_DATA_TEMPR67[22] , 
        \R_DATA_TEMPR67[21] , \R_DATA_TEMPR67[20] }), .B_DOUT({
        \R_DATA_TEMPR67[19] , \R_DATA_TEMPR67[18] , 
        \R_DATA_TEMPR67[17] , \R_DATA_TEMPR67[16] , 
        \R_DATA_TEMPR67[15] , \R_DATA_TEMPR67[14] , 
        \R_DATA_TEMPR67[13] , \R_DATA_TEMPR67[12] , 
        \R_DATA_TEMPR67[11] , \R_DATA_TEMPR67[10] , 
        \R_DATA_TEMPR67[9] , \R_DATA_TEMPR67[8] , \R_DATA_TEMPR67[7] , 
        \R_DATA_TEMPR67[6] , \R_DATA_TEMPR67[5] , \R_DATA_TEMPR67[4] , 
        \R_DATA_TEMPR67[3] , \R_DATA_TEMPR67[2] , \R_DATA_TEMPR67[1] , 
        \R_DATA_TEMPR67[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[67][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[16] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[16] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_622 (.A(\R_DATA_TEMPR96[5] ), .B(\R_DATA_TEMPR97[5] ), .C(
        \R_DATA_TEMPR98[5] ), .D(\R_DATA_TEMPR99[5] ), .Y(OR4_622_Y));
    OR4 OR4_232 (.A(\R_DATA_TEMPR108[2] ), .B(\R_DATA_TEMPR109[2] ), 
        .C(\R_DATA_TEMPR110[2] ), .D(\R_DATA_TEMPR111[2] ), .Y(
        OR4_232_Y));
    OR4 OR4_1579 (.A(OR4_666_Y), .B(OR4_501_Y), .C(OR4_1525_Y), .D(
        OR4_419_Y), .Y(OR4_1579_Y));
    OR4 OR4_844 (.A(\R_DATA_TEMPR64[29] ), .B(\R_DATA_TEMPR65[29] ), 
        .C(\R_DATA_TEMPR66[29] ), .D(\R_DATA_TEMPR67[29] ), .Y(
        OR4_844_Y));
    CFG3 #( .INIT(8'h2) )  CFG3_6 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_6_Y));
    OR4 \OR4_R_DATA[15]  (.A(OR4_1435_Y), .B(OR4_576_Y), .C(OR4_1196_Y)
        , .D(OR4_738_Y), .Y(R_DATA[15]));
    OR4 OR4_1167 (.A(OR4_726_Y), .B(OR4_1506_Y), .C(OR4_352_Y), .D(
        OR4_648_Y), .Y(OR4_1167_Y));
    OR4 OR4_543 (.A(\R_DATA_TEMPR116[21] ), .B(\R_DATA_TEMPR117[21] ), 
        .C(\R_DATA_TEMPR118[21] ), .D(\R_DATA_TEMPR119[21] ), .Y(
        OR4_543_Y));
    OR2 OR2_12 (.A(\R_DATA_TEMPR84[37] ), .B(\R_DATA_TEMPR85[37] ), .Y(
        OR2_12_Y));
    OR4 OR4_45 (.A(\R_DATA_TEMPR96[1] ), .B(\R_DATA_TEMPR97[1] ), .C(
        \R_DATA_TEMPR98[1] ), .D(\R_DATA_TEMPR99[1] ), .Y(OR4_45_Y));
    OR4 OR4_367 (.A(\R_DATA_TEMPR124[4] ), .B(\R_DATA_TEMPR125[4] ), 
        .C(\R_DATA_TEMPR126[4] ), .D(\R_DATA_TEMPR127[4] ), .Y(
        OR4_367_Y));
    OR4 OR4_160 (.A(\R_DATA_TEMPR12[21] ), .B(\R_DATA_TEMPR13[21] ), 
        .C(\R_DATA_TEMPR14[21] ), .D(\R_DATA_TEMPR15[21] ), .Y(
        OR4_160_Y));
    OR4 OR4_702 (.A(OR4_67_Y), .B(OR4_1520_Y), .C(OR4_914_Y), .D(
        OR4_1454_Y), .Y(OR4_702_Y));
    OR4 OR4_559 (.A(\R_DATA_TEMPR72[26] ), .B(\R_DATA_TEMPR73[26] ), 
        .C(\R_DATA_TEMPR74[26] ), .D(\R_DATA_TEMPR75[26] ), .Y(
        OR4_559_Y));
    OR4 OR4_1044 (.A(\R_DATA_TEMPR100[37] ), .B(\R_DATA_TEMPR101[37] ), 
        .C(\R_DATA_TEMPR102[37] ), .D(\R_DATA_TEMPR103[37] ), .Y(
        OR4_1044_Y));
    OR4 OR4_550 (.A(\R_DATA_TEMPR108[34] ), .B(\R_DATA_TEMPR109[34] ), 
        .C(\R_DATA_TEMPR110[34] ), .D(\R_DATA_TEMPR111[34] ), .Y(
        OR4_550_Y));
    OR4 \OR4_R_DATA[23]  (.A(OR4_865_Y), .B(OR4_441_Y), .C(OR4_375_Y), 
        .D(OR4_335_Y), .Y(R_DATA[23]));
    OR4 OR4_1583 (.A(\R_DATA_TEMPR12[28] ), .B(\R_DATA_TEMPR13[28] ), 
        .C(\R_DATA_TEMPR14[28] ), .D(\R_DATA_TEMPR15[28] ), .Y(
        OR4_1583_Y));
    OR4 OR4_330 (.A(OR4_123_Y), .B(OR4_1287_Y), .C(OR4_187_Y), .D(
        OR4_642_Y), .Y(OR4_330_Y));
    OR4 OR4_906 (.A(OR4_762_Y), .B(OR2_2_Y), .C(\R_DATA_TEMPR86[25] ), 
        .D(\R_DATA_TEMPR87[25] ), .Y(OR4_906_Y));
    OR4 OR4_772 (.A(OR4_849_Y), .B(OR4_1433_Y), .C(OR4_583_Y), .D(
        OR4_832_Y), .Y(OR4_772_Y));
    OR4 OR4_768 (.A(\R_DATA_TEMPR76[12] ), .B(\R_DATA_TEMPR77[12] ), 
        .C(\R_DATA_TEMPR78[12] ), .D(\R_DATA_TEMPR79[12] ), .Y(
        OR4_768_Y));
    OR4 OR4_1343 (.A(OR4_479_Y), .B(OR4_519_Y), .C(OR4_492_Y), .D(
        OR4_1265_Y), .Y(OR4_1343_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%16%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C0 (.A_DOUT({
        \R_DATA_TEMPR16[39] , \R_DATA_TEMPR16[38] , 
        \R_DATA_TEMPR16[37] , \R_DATA_TEMPR16[36] , 
        \R_DATA_TEMPR16[35] , \R_DATA_TEMPR16[34] , 
        \R_DATA_TEMPR16[33] , \R_DATA_TEMPR16[32] , 
        \R_DATA_TEMPR16[31] , \R_DATA_TEMPR16[30] , 
        \R_DATA_TEMPR16[29] , \R_DATA_TEMPR16[28] , 
        \R_DATA_TEMPR16[27] , \R_DATA_TEMPR16[26] , 
        \R_DATA_TEMPR16[25] , \R_DATA_TEMPR16[24] , 
        \R_DATA_TEMPR16[23] , \R_DATA_TEMPR16[22] , 
        \R_DATA_TEMPR16[21] , \R_DATA_TEMPR16[20] }), .B_DOUT({
        \R_DATA_TEMPR16[19] , \R_DATA_TEMPR16[18] , 
        \R_DATA_TEMPR16[17] , \R_DATA_TEMPR16[16] , 
        \R_DATA_TEMPR16[15] , \R_DATA_TEMPR16[14] , 
        \R_DATA_TEMPR16[13] , \R_DATA_TEMPR16[12] , 
        \R_DATA_TEMPR16[11] , \R_DATA_TEMPR16[10] , 
        \R_DATA_TEMPR16[9] , \R_DATA_TEMPR16[8] , \R_DATA_TEMPR16[7] , 
        \R_DATA_TEMPR16[6] , \R_DATA_TEMPR16[5] , \R_DATA_TEMPR16[4] , 
        \R_DATA_TEMPR16[3] , \R_DATA_TEMPR16[2] , \R_DATA_TEMPR16[1] , 
        \R_DATA_TEMPR16[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_605 (.A(OR4_586_Y), .B(OR4_333_Y), .C(OR4_31_Y), .D(
        OR4_50_Y), .Y(OR4_605_Y));
    OR4 OR4_511 (.A(\R_DATA_TEMPR124[38] ), .B(\R_DATA_TEMPR125[38] ), 
        .C(\R_DATA_TEMPR126[38] ), .D(\R_DATA_TEMPR127[38] ), .Y(
        OR4_511_Y));
    OR4 OR4_976 (.A(\R_DATA_TEMPR76[16] ), .B(\R_DATA_TEMPR77[16] ), 
        .C(\R_DATA_TEMPR78[16] ), .D(\R_DATA_TEMPR79[16] ), .Y(
        OR4_976_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[20]  (.A(CFG3_6_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[20] ));
    OR4 OR4_1415 (.A(OR4_683_Y), .B(OR4_530_Y), .C(OR4_649_Y), .D(
        OR4_751_Y), .Y(OR4_1415_Y));
    OR4 OR4_1233 (.A(\R_DATA_TEMPR56[13] ), .B(\R_DATA_TEMPR57[13] ), 
        .C(\R_DATA_TEMPR58[13] ), .D(\R_DATA_TEMPR59[13] ), .Y(
        OR4_1233_Y));
    OR4 OR4_833 (.A(\R_DATA_TEMPR72[28] ), .B(\R_DATA_TEMPR73[28] ), 
        .C(\R_DATA_TEMPR74[28] ), .D(\R_DATA_TEMPR75[28] ), .Y(
        OR4_833_Y));
    OR4 OR4_825 (.A(\R_DATA_TEMPR52[28] ), .B(\R_DATA_TEMPR53[28] ), 
        .C(\R_DATA_TEMPR54[28] ), .D(\R_DATA_TEMPR55[28] ), .Y(
        OR4_825_Y));
    OR4 OR4_696 (.A(\R_DATA_TEMPR20[30] ), .B(\R_DATA_TEMPR21[30] ), 
        .C(\R_DATA_TEMPR22[30] ), .D(\R_DATA_TEMPR23[30] ), .Y(
        OR4_696_Y));
    OR4 OR4_675 (.A(OR4_993_Y), .B(OR4_1581_Y), .C(OR4_729_Y), .D(
        OR4_984_Y), .Y(OR4_675_Y));
    OR4 OR4_287 (.A(\R_DATA_TEMPR4[13] ), .B(\R_DATA_TEMPR5[13] ), .C(
        \R_DATA_TEMPR6[13] ), .D(\R_DATA_TEMPR7[13] ), .Y(OR4_287_Y));
    OR4 OR4_86 (.A(\R_DATA_TEMPR116[1] ), .B(\R_DATA_TEMPR117[1] ), .C(
        \R_DATA_TEMPR118[1] ), .D(\R_DATA_TEMPR119[1] ), .Y(OR4_86_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[4]  (.A(CFG3_6_Y), .B(CFG3_12_Y)
        , .Y(\BLKX2[4] ));
    OR4 OR4_33 (.A(OR4_1449_Y), .B(OR4_109_Y), .C(OR4_1188_Y), .D(
        OR4_422_Y), .Y(OR4_33_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[10]  (.A(CFG3_0_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[10] ));
    OR4 OR4_867 (.A(\R_DATA_TEMPR120[32] ), .B(\R_DATA_TEMPR121[32] ), 
        .C(\R_DATA_TEMPR122[32] ), .D(\R_DATA_TEMPR123[32] ), .Y(
        OR4_867_Y));
    OR4 OR4_168 (.A(\R_DATA_TEMPR108[32] ), .B(\R_DATA_TEMPR109[32] ), 
        .C(\R_DATA_TEMPR110[32] ), .D(\R_DATA_TEMPR111[32] ), .Y(
        OR4_168_Y));
    OR4 OR4_964 (.A(\R_DATA_TEMPR116[30] ), .B(\R_DATA_TEMPR117[30] ), 
        .C(\R_DATA_TEMPR118[30] ), .D(\R_DATA_TEMPR119[30] ), .Y(
        OR4_964_Y));
    OR4 OR4_187 (.A(\R_DATA_TEMPR88[4] ), .B(\R_DATA_TEMPR89[4] ), .C(
        \R_DATA_TEMPR90[4] ), .D(\R_DATA_TEMPR91[4] ), .Y(OR4_187_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%97%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R97C0 (.A_DOUT({
        \R_DATA_TEMPR97[39] , \R_DATA_TEMPR97[38] , 
        \R_DATA_TEMPR97[37] , \R_DATA_TEMPR97[36] , 
        \R_DATA_TEMPR97[35] , \R_DATA_TEMPR97[34] , 
        \R_DATA_TEMPR97[33] , \R_DATA_TEMPR97[32] , 
        \R_DATA_TEMPR97[31] , \R_DATA_TEMPR97[30] , 
        \R_DATA_TEMPR97[29] , \R_DATA_TEMPR97[28] , 
        \R_DATA_TEMPR97[27] , \R_DATA_TEMPR97[26] , 
        \R_DATA_TEMPR97[25] , \R_DATA_TEMPR97[24] , 
        \R_DATA_TEMPR97[23] , \R_DATA_TEMPR97[22] , 
        \R_DATA_TEMPR97[21] , \R_DATA_TEMPR97[20] }), .B_DOUT({
        \R_DATA_TEMPR97[19] , \R_DATA_TEMPR97[18] , 
        \R_DATA_TEMPR97[17] , \R_DATA_TEMPR97[16] , 
        \R_DATA_TEMPR97[15] , \R_DATA_TEMPR97[14] , 
        \R_DATA_TEMPR97[13] , \R_DATA_TEMPR97[12] , 
        \R_DATA_TEMPR97[11] , \R_DATA_TEMPR97[10] , 
        \R_DATA_TEMPR97[9] , \R_DATA_TEMPR97[8] , \R_DATA_TEMPR97[7] , 
        \R_DATA_TEMPR97[6] , \R_DATA_TEMPR97[5] , \R_DATA_TEMPR97[4] , 
        \R_DATA_TEMPR97[3] , \R_DATA_TEMPR97[2] , \R_DATA_TEMPR97[1] , 
        \R_DATA_TEMPR97[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[97][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[24] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[24] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1052 (.A(\R_DATA_TEMPR92[21] ), .B(\R_DATA_TEMPR93[21] ), 
        .C(\R_DATA_TEMPR94[21] ), .D(\R_DATA_TEMPR95[21] ), .Y(
        OR4_1052_Y));
    OR4 OR4_212 (.A(\R_DATA_TEMPR92[8] ), .B(\R_DATA_TEMPR93[8] ), .C(
        \R_DATA_TEMPR94[8] ), .D(\R_DATA_TEMPR95[8] ), .Y(OR4_212_Y));
    OR4 OR4_1197 (.A(\R_DATA_TEMPR8[3] ), .B(\R_DATA_TEMPR9[3] ), .C(
        \R_DATA_TEMPR10[3] ), .D(\R_DATA_TEMPR11[3] ), .Y(OR4_1197_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%9%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C0 (.A_DOUT({
        \R_DATA_TEMPR9[39] , \R_DATA_TEMPR9[38] , \R_DATA_TEMPR9[37] , 
        \R_DATA_TEMPR9[36] , \R_DATA_TEMPR9[35] , \R_DATA_TEMPR9[34] , 
        \R_DATA_TEMPR9[33] , \R_DATA_TEMPR9[32] , \R_DATA_TEMPR9[31] , 
        \R_DATA_TEMPR9[30] , \R_DATA_TEMPR9[29] , \R_DATA_TEMPR9[28] , 
        \R_DATA_TEMPR9[27] , \R_DATA_TEMPR9[26] , \R_DATA_TEMPR9[25] , 
        \R_DATA_TEMPR9[24] , \R_DATA_TEMPR9[23] , \R_DATA_TEMPR9[22] , 
        \R_DATA_TEMPR9[21] , \R_DATA_TEMPR9[20] }), .B_DOUT({
        \R_DATA_TEMPR9[19] , \R_DATA_TEMPR9[18] , \R_DATA_TEMPR9[17] , 
        \R_DATA_TEMPR9[16] , \R_DATA_TEMPR9[15] , \R_DATA_TEMPR9[14] , 
        \R_DATA_TEMPR9[13] , \R_DATA_TEMPR9[12] , \R_DATA_TEMPR9[11] , 
        \R_DATA_TEMPR9[10] , \R_DATA_TEMPR9[9] , \R_DATA_TEMPR9[8] , 
        \R_DATA_TEMPR9[7] , \R_DATA_TEMPR9[6] , \R_DATA_TEMPR9[5] , 
        \R_DATA_TEMPR9[4] , \R_DATA_TEMPR9[3] , \R_DATA_TEMPR9[2] , 
        \R_DATA_TEMPR9[1] , \R_DATA_TEMPR9[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[9][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1575 (.A(\R_DATA_TEMPR124[14] ), .B(\R_DATA_TEMPR125[14] ), 
        .C(\R_DATA_TEMPR126[14] ), .D(\R_DATA_TEMPR127[14] ), .Y(
        OR4_1575_Y));
    OR4 OR4_1614 (.A(\R_DATA_TEMPR52[9] ), .B(\R_DATA_TEMPR53[9] ), .C(
        \R_DATA_TEMPR54[9] ), .D(\R_DATA_TEMPR55[9] ), .Y(OR4_1614_Y));
    OR4 OR4_353 (.A(\R_DATA_TEMPR76[24] ), .B(\R_DATA_TEMPR77[24] ), 
        .C(\R_DATA_TEMPR78[24] ), .D(\R_DATA_TEMPR79[24] ), .Y(
        OR4_353_Y));
    OR4 OR4_1139 (.A(OR4_132_Y), .B(OR4_900_Y), .C(OR4_871_Y), .D(
        OR4_9_Y), .Y(OR4_1139_Y));
    OR4 OR4_750 (.A(\R_DATA_TEMPR52[23] ), .B(\R_DATA_TEMPR53[23] ), 
        .C(\R_DATA_TEMPR54[23] ), .D(\R_DATA_TEMPR55[23] ), .Y(
        OR4_750_Y));
    OR4 OR4_1260 (.A(\R_DATA_TEMPR32[17] ), .B(\R_DATA_TEMPR33[17] ), 
        .C(\R_DATA_TEMPR34[17] ), .D(\R_DATA_TEMPR35[17] ), .Y(
        OR4_1260_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[2]  (.A(CFG3_0_Y), .B(CFG3_2_Y), 
        .Y(\BLKY2[2] ));
    OR4 OR4_783 (.A(\R_DATA_TEMPR88[26] ), .B(\R_DATA_TEMPR89[26] ), 
        .C(\R_DATA_TEMPR90[26] ), .D(\R_DATA_TEMPR91[26] ), .Y(
        OR4_783_Y));
    OR4 OR4_1276 (.A(\R_DATA_TEMPR28[36] ), .B(\R_DATA_TEMPR29[36] ), 
        .C(\R_DATA_TEMPR30[36] ), .D(\R_DATA_TEMPR31[36] ), .Y(
        OR4_1276_Y));
    OR4 OR4_600 (.A(\R_DATA_TEMPR68[18] ), .B(\R_DATA_TEMPR69[18] ), 
        .C(\R_DATA_TEMPR70[18] ), .D(\R_DATA_TEMPR71[18] ), .Y(
        OR4_600_Y));
    OR4 OR4_452 (.A(\R_DATA_TEMPR60[17] ), .B(\R_DATA_TEMPR61[17] ), 
        .C(\R_DATA_TEMPR62[17] ), .D(\R_DATA_TEMPR63[17] ), .Y(
        OR4_452_Y));
    OR4 OR4_284 (.A(OR4_673_Y), .B(OR4_518_Y), .C(OR4_639_Y), .D(
        OR4_1039_Y), .Y(OR4_284_Y));
    OR4 OR4_310 (.A(OR4_28_Y), .B(OR4_378_Y), .C(OR4_561_Y), .D(
        OR4_113_Y), .Y(OR4_310_Y));
    OR4 OR4_5 (.A(\R_DATA_TEMPR16[1] ), .B(\R_DATA_TEMPR17[1] ), .C(
        \R_DATA_TEMPR18[1] ), .D(\R_DATA_TEMPR19[1] ), .Y(OR4_5_Y));
    OR4 OR4_1316 (.A(\R_DATA_TEMPR8[17] ), .B(\R_DATA_TEMPR9[17] ), .C(
        \R_DATA_TEMPR10[17] ), .D(\R_DATA_TEMPR11[17] ), .Y(OR4_1316_Y)
        );
    OR4 OR4_1403 (.A(\R_DATA_TEMPR88[8] ), .B(\R_DATA_TEMPR89[8] ), .C(
        \R_DATA_TEMPR90[8] ), .D(\R_DATA_TEMPR91[8] ), .Y(OR4_1403_Y));
    OR4 OR4_1378 (.A(\R_DATA_TEMPR8[20] ), .B(\R_DATA_TEMPR9[20] ), .C(
        \R_DATA_TEMPR10[20] ), .D(\R_DATA_TEMPR11[20] ), .Y(OR4_1378_Y)
        );
    OR4 OR4_1046 (.A(\R_DATA_TEMPR108[19] ), .B(\R_DATA_TEMPR109[19] ), 
        .C(\R_DATA_TEMPR110[19] ), .D(\R_DATA_TEMPR111[19] ), .Y(
        OR4_1046_Y));
    OR4 OR4_670 (.A(OR4_539_Y), .B(OR4_785_Y), .C(OR4_304_Y), .D(
        OR4_29_Y), .Y(OR4_670_Y));
    OR4 OR4_1567 (.A(\R_DATA_TEMPR124[1] ), .B(\R_DATA_TEMPR125[1] ), 
        .C(\R_DATA_TEMPR126[1] ), .D(\R_DATA_TEMPR127[1] ), .Y(
        OR4_1567_Y));
    OR4 OR4_459 (.A(\R_DATA_TEMPR116[24] ), .B(\R_DATA_TEMPR117[24] ), 
        .C(\R_DATA_TEMPR118[24] ), .D(\R_DATA_TEMPR119[24] ), .Y(
        OR4_459_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[27]  (.A(CFG3_19_Y), .B(
        CFG3_3_Y), .Y(\BLKY2[27] ));
    OR4 OR4_307 (.A(\R_DATA_TEMPR56[15] ), .B(\R_DATA_TEMPR57[15] ), 
        .C(\R_DATA_TEMPR58[15] ), .D(\R_DATA_TEMPR59[15] ), .Y(
        OR4_307_Y));
    OR4 OR4_100 (.A(\R_DATA_TEMPR36[6] ), .B(\R_DATA_TEMPR37[6] ), .C(
        \R_DATA_TEMPR38[6] ), .D(\R_DATA_TEMPR39[6] ), .Y(OR4_100_Y));
    OR4 OR4_1611 (.A(\R_DATA_TEMPR72[0] ), .B(\R_DATA_TEMPR73[0] ), .C(
        \R_DATA_TEMPR74[0] ), .D(\R_DATA_TEMPR75[0] ), .Y(OR4_1611_Y));
    OR4 OR4_1362 (.A(OR4_150_Y), .B(OR4_713_Y), .C(OR4_690_Y), .D(
        OR4_376_Y), .Y(OR4_1362_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[28]  (.A(CFG3_6_Y), .B(CFG3_7_Y)
        , .Y(\BLKX2[28] ));
    OR4 OR4_99 (.A(\R_DATA_TEMPR24[11] ), .B(\R_DATA_TEMPR25[11] ), .C(
        \R_DATA_TEMPR26[11] ), .D(\R_DATA_TEMPR27[11] ), .Y(OR4_99_Y));
    OR4 OR4_156 (.A(\R_DATA_TEMPR100[28] ), .B(\R_DATA_TEMPR101[28] ), 
        .C(\R_DATA_TEMPR102[28] ), .D(\R_DATA_TEMPR103[28] ), .Y(
        OR4_156_Y));
    OR4 OR4_1223 (.A(\R_DATA_TEMPR100[39] ), .B(\R_DATA_TEMPR101[39] ), 
        .C(\R_DATA_TEMPR102[39] ), .D(\R_DATA_TEMPR103[39] ), .Y(
        OR4_1223_Y));
    OR4 OR4_535 (.A(\R_DATA_TEMPR112[3] ), .B(\R_DATA_TEMPR113[3] ), 
        .C(\R_DATA_TEMPR114[3] ), .D(\R_DATA_TEMPR115[3] ), .Y(
        OR4_535_Y));
    OR2 OR2_36 (.A(\R_DATA_TEMPR84[23] ), .B(\R_DATA_TEMPR85[23] ), .Y(
        OR2_36_Y));
    OR4 OR4_1262 (.A(\R_DATA_TEMPR24[32] ), .B(\R_DATA_TEMPR25[32] ), 
        .C(\R_DATA_TEMPR26[32] ), .D(\R_DATA_TEMPR27[32] ), .Y(
        OR4_1262_Y));
    OR4 OR4_813 (.A(OR4_1511_Y), .B(OR4_189_Y), .C(OR4_433_Y), .D(
        OR4_240_Y), .Y(OR4_813_Y));
    OR2 OR2_24 (.A(\R_DATA_TEMPR84[36] ), .B(\R_DATA_TEMPR85[36] ), .Y(
        OR2_24_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[23]  (.A(CFG3_23_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[23] ));
    OR4 OR4_68 (.A(\R_DATA_TEMPR64[22] ), .B(\R_DATA_TEMPR65[22] ), .C(
        \R_DATA_TEMPR66[22] ), .D(\R_DATA_TEMPR67[22] ), .Y(OR4_68_Y));
    OR4 OR4_377 (.A(\R_DATA_TEMPR16[24] ), .B(\R_DATA_TEMPR17[24] ), 
        .C(\R_DATA_TEMPR18[24] ), .D(\R_DATA_TEMPR19[24] ), .Y(
        OR4_377_Y));
    OR4 OR4_170 (.A(OR4_1355_Y), .B(OR4_1173_Y), .C(OR4_1324_Y), .D(
        OR4_98_Y), .Y(OR4_170_Y));
    OR4 OR4_1610 (.A(\R_DATA_TEMPR64[20] ), .B(\R_DATA_TEMPR65[20] ), 
        .C(\R_DATA_TEMPR66[20] ), .D(\R_DATA_TEMPR67[20] ), .Y(
        OR4_1610_Y));
    OR4 OR4_1341 (.A(\R_DATA_TEMPR28[30] ), .B(\R_DATA_TEMPR29[30] ), 
        .C(\R_DATA_TEMPR30[30] ), .D(\R_DATA_TEMPR31[30] ), .Y(
        OR4_1341_Y));
    OR4 OR4_708 (.A(\R_DATA_TEMPR36[37] ), .B(\R_DATA_TEMPR37[37] ), 
        .C(\R_DATA_TEMPR38[37] ), .D(\R_DATA_TEMPR39[37] ), .Y(
        OR4_708_Y));
    OR4 OR4_626 (.A(\R_DATA_TEMPR100[38] ), .B(\R_DATA_TEMPR101[38] ), 
        .C(\R_DATA_TEMPR102[38] ), .D(\R_DATA_TEMPR103[38] ), .Y(
        OR4_626_Y));
    OR4 OR4_31 (.A(\R_DATA_TEMPR120[25] ), .B(\R_DATA_TEMPR121[25] ), 
        .C(\R_DATA_TEMPR122[25] ), .D(\R_DATA_TEMPR123[25] ), .Y(
        OR4_31_Y));
    OR4 OR4_633 (.A(\R_DATA_TEMPR16[9] ), .B(\R_DATA_TEMPR17[9] ), .C(
        \R_DATA_TEMPR18[9] ), .D(\R_DATA_TEMPR19[9] ), .Y(OR4_633_Y));
    OR4 OR4_1464 (.A(\R_DATA_TEMPR76[14] ), .B(\R_DATA_TEMPR77[14] ), 
        .C(\R_DATA_TEMPR78[14] ), .D(\R_DATA_TEMPR79[14] ), .Y(
        OR4_1464_Y));
    OR4 \OR4_R_DATA[31]  (.A(OR4_389_Y), .B(OR4_319_Y), .C(OR4_342_Y), 
        .D(OR4_1470_Y), .Y(R_DATA[31]));
    OR4 OR4_1136 (.A(\R_DATA_TEMPR52[22] ), .B(\R_DATA_TEMPR53[22] ), 
        .C(\R_DATA_TEMPR54[22] ), .D(\R_DATA_TEMPR55[22] ), .Y(
        OR4_1136_Y));
    OR4 OR4_385 (.A(\R_DATA_TEMPR4[31] ), .B(\R_DATA_TEMPR5[31] ), .C(
        \R_DATA_TEMPR6[31] ), .D(\R_DATA_TEMPR7[31] ), .Y(OR4_385_Y));
    OR4 OR4_778 (.A(\R_DATA_TEMPR12[30] ), .B(\R_DATA_TEMPR13[30] ), 
        .C(\R_DATA_TEMPR14[30] ), .D(\R_DATA_TEMPR15[30] ), .Y(
        OR4_778_Y));
    OR4 OR4_1431 (.A(OR4_917_Y), .B(OR4_587_Y), .C(OR4_326_Y), .D(
        OR4_394_Y), .Y(OR4_1431_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[15]  (.A(CFG3_23_Y), .B(
        CFG3_4_Y), .Y(\BLKX2[15] ));
    OR4 OR4_243 (.A(\R_DATA_TEMPR76[31] ), .B(\R_DATA_TEMPR77[31] ), 
        .C(\R_DATA_TEMPR78[31] ), .D(\R_DATA_TEMPR79[31] ), .Y(
        OR4_243_Y));
    OR4 OR4_394 (.A(OR4_260_Y), .B(OR4_825_Y), .C(OR4_1622_Y), .D(
        OR4_244_Y), .Y(OR4_394_Y));
    OR4 OR4_1079 (.A(\R_DATA_TEMPR36[7] ), .B(\R_DATA_TEMPR37[7] ), .C(
        \R_DATA_TEMPR38[7] ), .D(\R_DATA_TEMPR39[7] ), .Y(OR4_1079_Y));
    OR4 OR4_1264 (.A(\R_DATA_TEMPR32[12] ), .B(\R_DATA_TEMPR33[12] ), 
        .C(\R_DATA_TEMPR34[12] ), .D(\R_DATA_TEMPR35[12] ), .Y(
        OR4_1264_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%36%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R36C0 (.A_DOUT({
        \R_DATA_TEMPR36[39] , \R_DATA_TEMPR36[38] , 
        \R_DATA_TEMPR36[37] , \R_DATA_TEMPR36[36] , 
        \R_DATA_TEMPR36[35] , \R_DATA_TEMPR36[34] , 
        \R_DATA_TEMPR36[33] , \R_DATA_TEMPR36[32] , 
        \R_DATA_TEMPR36[31] , \R_DATA_TEMPR36[30] , 
        \R_DATA_TEMPR36[29] , \R_DATA_TEMPR36[28] , 
        \R_DATA_TEMPR36[27] , \R_DATA_TEMPR36[26] , 
        \R_DATA_TEMPR36[25] , \R_DATA_TEMPR36[24] , 
        \R_DATA_TEMPR36[23] , \R_DATA_TEMPR36[22] , 
        \R_DATA_TEMPR36[21] , \R_DATA_TEMPR36[20] }), .B_DOUT({
        \R_DATA_TEMPR36[19] , \R_DATA_TEMPR36[18] , 
        \R_DATA_TEMPR36[17] , \R_DATA_TEMPR36[16] , 
        \R_DATA_TEMPR36[15] , \R_DATA_TEMPR36[14] , 
        \R_DATA_TEMPR36[13] , \R_DATA_TEMPR36[12] , 
        \R_DATA_TEMPR36[11] , \R_DATA_TEMPR36[10] , 
        \R_DATA_TEMPR36[9] , \R_DATA_TEMPR36[8] , \R_DATA_TEMPR36[7] , 
        \R_DATA_TEMPR36[6] , \R_DATA_TEMPR36[5] , \R_DATA_TEMPR36[4] , 
        \R_DATA_TEMPR36[3] , \R_DATA_TEMPR36[2] , \R_DATA_TEMPR36[1] , 
        \R_DATA_TEMPR36[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[36][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[9] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[9] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_358 (.A(OR4_1143_Y), .B(OR4_558_Y), .C(OR4_791_Y), .D(
        OR4_1380_Y), .Y(OR4_358_Y));
    OR4 OR4_1483 (.A(\R_DATA_TEMPR32[18] ), .B(\R_DATA_TEMPR33[18] ), 
        .C(\R_DATA_TEMPR34[18] ), .D(\R_DATA_TEMPR35[18] ), .Y(
        OR4_1483_Y));
    OR4 OR4_1231 (.A(\R_DATA_TEMPR16[37] ), .B(\R_DATA_TEMPR17[37] ), 
        .C(\R_DATA_TEMPR18[37] ), .D(\R_DATA_TEMPR19[37] ), .Y(
        OR4_1231_Y));
    OR4 OR4_1553 (.A(OR4_267_Y), .B(OR4_321_Y), .C(OR4_836_Y), .D(
        OR4_1289_Y), .Y(OR4_1553_Y));
    OR4 OR4_1138 (.A(OR4_1264_Y), .B(OR4_1501_Y), .C(OR4_1479_Y), .D(
        OR4_616_Y), .Y(OR4_1138_Y));
    OR4 OR4_80 (.A(\R_DATA_TEMPR16[14] ), .B(\R_DATA_TEMPR17[14] ), .C(
        \R_DATA_TEMPR18[14] ), .D(\R_DATA_TEMPR19[14] ), .Y(OR4_80_Y));
    OR4 OR4_1367 (.A(\R_DATA_TEMPR108[3] ), .B(\R_DATA_TEMPR109[3] ), 
        .C(\R_DATA_TEMPR110[3] ), .D(\R_DATA_TEMPR111[3] ), .Y(
        OR4_1367_Y));
    OR4 OR4_807 (.A(\R_DATA_TEMPR124[36] ), .B(\R_DATA_TEMPR125[36] ), 
        .C(\R_DATA_TEMPR126[36] ), .D(\R_DATA_TEMPR127[36] ), .Y(
        OR4_807_Y));
    OR4 OR4_108 (.A(\R_DATA_TEMPR44[3] ), .B(\R_DATA_TEMPR45[3] ), .C(
        \R_DATA_TEMPR46[3] ), .D(\R_DATA_TEMPR47[3] ), .Y(OR4_108_Y));
    OR4 OR4_191 (.A(\R_DATA_TEMPR64[6] ), .B(\R_DATA_TEMPR65[6] ), .C(
        \R_DATA_TEMPR66[6] ), .D(\R_DATA_TEMPR67[6] ), .Y(OR4_191_Y));
    OR4 OR4_1290 (.A(\R_DATA_TEMPR76[22] ), .B(\R_DATA_TEMPR77[22] ), 
        .C(\R_DATA_TEMPR78[22] ), .D(\R_DATA_TEMPR79[22] ), .Y(
        OR4_1290_Y));
    OR4 OR4_1129 (.A(\R_DATA_TEMPR112[27] ), .B(\R_DATA_TEMPR113[27] ), 
        .C(\R_DATA_TEMPR114[27] ), .D(\R_DATA_TEMPR115[27] ), .Y(
        OR4_1129_Y));
    OR4 OR4_904 (.A(OR4_1486_Y), .B(OR4_1301_Y), .C(OR4_688_Y), .D(
        OR4_1213_Y), .Y(OR4_904_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%69%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R69C0 (.A_DOUT({
        \R_DATA_TEMPR69[39] , \R_DATA_TEMPR69[38] , 
        \R_DATA_TEMPR69[37] , \R_DATA_TEMPR69[36] , 
        \R_DATA_TEMPR69[35] , \R_DATA_TEMPR69[34] , 
        \R_DATA_TEMPR69[33] , \R_DATA_TEMPR69[32] , 
        \R_DATA_TEMPR69[31] , \R_DATA_TEMPR69[30] , 
        \R_DATA_TEMPR69[29] , \R_DATA_TEMPR69[28] , 
        \R_DATA_TEMPR69[27] , \R_DATA_TEMPR69[26] , 
        \R_DATA_TEMPR69[25] , \R_DATA_TEMPR69[24] , 
        \R_DATA_TEMPR69[23] , \R_DATA_TEMPR69[22] , 
        \R_DATA_TEMPR69[21] , \R_DATA_TEMPR69[20] }), .B_DOUT({
        \R_DATA_TEMPR69[19] , \R_DATA_TEMPR69[18] , 
        \R_DATA_TEMPR69[17] , \R_DATA_TEMPR69[16] , 
        \R_DATA_TEMPR69[15] , \R_DATA_TEMPR69[14] , 
        \R_DATA_TEMPR69[13] , \R_DATA_TEMPR69[12] , 
        \R_DATA_TEMPR69[11] , \R_DATA_TEMPR69[10] , 
        \R_DATA_TEMPR69[9] , \R_DATA_TEMPR69[8] , \R_DATA_TEMPR69[7] , 
        \R_DATA_TEMPR69[6] , \R_DATA_TEMPR69[5] , \R_DATA_TEMPR69[4] , 
        \R_DATA_TEMPR69[3] , \R_DATA_TEMPR69[2] , \R_DATA_TEMPR69[1] , 
        \R_DATA_TEMPR69[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[69][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[17] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[17] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1418 (.A(\R_DATA_TEMPR36[10] ), .B(\R_DATA_TEMPR37[10] ), 
        .C(\R_DATA_TEMPR38[10] ), .D(\R_DATA_TEMPR39[10] ), .Y(
        OR4_1418_Y));
    OR4 OR4_948 (.A(\R_DATA_TEMPR112[8] ), .B(\R_DATA_TEMPR113[8] ), 
        .C(\R_DATA_TEMPR114[8] ), .D(\R_DATA_TEMPR115[8] ), .Y(
        OR4_948_Y));
    OR4 OR4_1 (.A(\R_DATA_TEMPR44[28] ), .B(\R_DATA_TEMPR45[28] ), .C(
        \R_DATA_TEMPR46[28] ), .D(\R_DATA_TEMPR47[28] ), .Y(OR4_1_Y));
    OR4 OR4_87 (.A(\R_DATA_TEMPR72[11] ), .B(\R_DATA_TEMPR73[11] ), .C(
        \R_DATA_TEMPR74[11] ), .D(\R_DATA_TEMPR75[11] ), .Y(OR4_87_Y));
    OR4 \OR4_R_DATA[30]  (.A(OR4_84_Y), .B(OR4_454_Y), .C(OR4_1185_Y), 
        .D(OR4_572_Y), .Y(R_DATA[30]));
    OR4 OR4_877 (.A(OR4_1595_Y), .B(OR4_643_Y), .C(OR4_1168_Y), .D(
        OR4_1633_Y), .Y(OR4_877_Y));
    OR4 OR4_178 (.A(\R_DATA_TEMPR96[11] ), .B(\R_DATA_TEMPR97[11] ), 
        .C(\R_DATA_TEMPR98[11] ), .D(\R_DATA_TEMPR99[11] ), .Y(
        OR4_178_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[0]  (.A(CFG3_13_Y), .B(
        CFG3_12_Y), .Y(\BLKX2[0] ));
    OR4 OR4_974 (.A(\R_DATA_TEMPR24[3] ), .B(\R_DATA_TEMPR25[3] ), .C(
        \R_DATA_TEMPR26[3] ), .D(\R_DATA_TEMPR27[3] ), .Y(OR4_974_Y));
    OR4 OR4_939 (.A(OR4_584_Y), .B(OR4_887_Y), .C(OR4_350_Y), .D(
        OR4_1182_Y), .Y(OR4_939_Y));
    OR4 OR4_930 (.A(\R_DATA_TEMPR96[16] ), .B(\R_DATA_TEMPR97[16] ), 
        .C(\R_DATA_TEMPR98[16] ), .D(\R_DATA_TEMPR99[16] ), .Y(
        OR4_930_Y));
    OR4 OR4_1597 (.A(\R_DATA_TEMPR60[26] ), .B(\R_DATA_TEMPR61[26] ), 
        .C(\R_DATA_TEMPR62[26] ), .D(\R_DATA_TEMPR63[26] ), .Y(
        OR4_1597_Y));
    OR4 OR4_1392 (.A(\R_DATA_TEMPR32[22] ), .B(\R_DATA_TEMPR33[22] ), 
        .C(\R_DATA_TEMPR34[22] ), .D(\R_DATA_TEMPR35[22] ), .Y(
        OR4_1392_Y));
    OR4 OR4_782 (.A(\R_DATA_TEMPR20[27] ), .B(\R_DATA_TEMPR21[27] ), 
        .C(\R_DATA_TEMPR22[27] ), .D(\R_DATA_TEMPR23[27] ), .Y(
        OR4_782_Y));
    OR4 OR4_159 (.A(\R_DATA_TEMPR120[24] ), .B(\R_DATA_TEMPR121[24] ), 
        .C(\R_DATA_TEMPR122[24] ), .D(\R_DATA_TEMPR123[24] ), .Y(
        OR4_159_Y));
    OR4 OR4_491 (.A(\R_DATA_TEMPR68[21] ), .B(\R_DATA_TEMPR69[21] ), 
        .C(\R_DATA_TEMPR70[21] ), .D(\R_DATA_TEMPR71[21] ), .Y(
        OR4_491_Y));
    OR4 OR4_165 (.A(\R_DATA_TEMPR32[21] ), .B(\R_DATA_TEMPR33[21] ), 
        .C(\R_DATA_TEMPR34[21] ), .D(\R_DATA_TEMPR35[21] ), .Y(
        OR4_165_Y));
    OR4 OR4_1292 (.A(OR4_487_Y), .B(OR4_927_Y), .C(OR4_271_Y), .D(
        OR4_580_Y), .Y(OR4_1292_Y));
    OR4 OR4_133 (.A(OR4_645_Y), .B(OR4_136_Y), .C(OR4_207_Y), .D(
        OR4_954_Y), .Y(OR4_133_Y));
    OR4 OR4_515 (.A(OR4_1160_Y), .B(OR4_1493_Y), .C(OR4_96_Y), .D(
        OR4_1531_Y), .Y(OR4_515_Y));
    OR4 OR4_498 (.A(\R_DATA_TEMPR100[11] ), .B(\R_DATA_TEMPR101[11] ), 
        .C(\R_DATA_TEMPR102[11] ), .D(\R_DATA_TEMPR103[11] ), .Y(
        OR4_498_Y));
    OR4 OR4_986 (.A(OR4_1389_Y), .B(OR2_4_Y), .C(\R_DATA_TEMPR86[7] ), 
        .D(\R_DATA_TEMPR87[7] ), .Y(OR4_986_Y));
    OR4 \OR4_R_DATA[36]  (.A(OR4_1131_Y), .B(OR4_397_Y), .C(OR4_676_Y), 
        .D(OR4_769_Y), .Y(R_DATA[36]));
    OR4 OR4_92 (.A(\R_DATA_TEMPR48[17] ), .B(\R_DATA_TEMPR49[17] ), .C(
        \R_DATA_TEMPR50[17] ), .D(\R_DATA_TEMPR51[17] ), .Y(OR4_92_Y));
    OR4 OR4_467 (.A(OR4_272_Y), .B(OR4_784_Y), .C(OR4_299_Y), .D(
        OR4_1439_Y), .Y(OR4_467_Y));
    OR4 OR4_1103 (.A(\R_DATA_TEMPR20[13] ), .B(\R_DATA_TEMPR21[13] ), 
        .C(\R_DATA_TEMPR22[13] ), .D(\R_DATA_TEMPR23[13] ), .Y(
        OR4_1103_Y));
    OR4 OR4_648 (.A(\R_DATA_TEMPR12[19] ), .B(\R_DATA_TEMPR13[19] ), 
        .C(\R_DATA_TEMPR14[19] ), .D(\R_DATA_TEMPR15[19] ), .Y(
        OR4_648_Y));
    OR4 OR4_1114 (.A(OR4_1098_Y), .B(OR2_11_Y), .C(
        \R_DATA_TEMPR86[21] ), .D(\R_DATA_TEMPR87[21] ), .Y(OR4_1114_Y)
        );
    OR4 OR4_685 (.A(\R_DATA_TEMPR96[19] ), .B(\R_DATA_TEMPR97[19] ), 
        .C(\R_DATA_TEMPR98[19] ), .D(\R_DATA_TEMPR99[19] ), .Y(
        OR4_685_Y));
    OR4 OR4_1494 (.A(\R_DATA_TEMPR112[0] ), .B(\R_DATA_TEMPR113[0] ), 
        .C(\R_DATA_TEMPR114[0] ), .D(\R_DATA_TEMPR115[0] ), .Y(
        OR4_1494_Y));
    OR4 OR4_613 (.A(\R_DATA_TEMPR40[28] ), .B(\R_DATA_TEMPR41[28] ), 
        .C(\R_DATA_TEMPR42[28] ), .D(\R_DATA_TEMPR43[28] ), .Y(
        OR4_613_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%104%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R104C0 (.A_DOUT({
        \R_DATA_TEMPR104[39] , \R_DATA_TEMPR104[38] , 
        \R_DATA_TEMPR104[37] , \R_DATA_TEMPR104[36] , 
        \R_DATA_TEMPR104[35] , \R_DATA_TEMPR104[34] , 
        \R_DATA_TEMPR104[33] , \R_DATA_TEMPR104[32] , 
        \R_DATA_TEMPR104[31] , \R_DATA_TEMPR104[30] , 
        \R_DATA_TEMPR104[29] , \R_DATA_TEMPR104[28] , 
        \R_DATA_TEMPR104[27] , \R_DATA_TEMPR104[26] , 
        \R_DATA_TEMPR104[25] , \R_DATA_TEMPR104[24] , 
        \R_DATA_TEMPR104[23] , \R_DATA_TEMPR104[22] , 
        \R_DATA_TEMPR104[21] , \R_DATA_TEMPR104[20] }), .B_DOUT({
        \R_DATA_TEMPR104[19] , \R_DATA_TEMPR104[18] , 
        \R_DATA_TEMPR104[17] , \R_DATA_TEMPR104[16] , 
        \R_DATA_TEMPR104[15] , \R_DATA_TEMPR104[14] , 
        \R_DATA_TEMPR104[13] , \R_DATA_TEMPR104[12] , 
        \R_DATA_TEMPR104[11] , \R_DATA_TEMPR104[10] , 
        \R_DATA_TEMPR104[9] , \R_DATA_TEMPR104[8] , 
        \R_DATA_TEMPR104[7] , \R_DATA_TEMPR104[6] , 
        \R_DATA_TEMPR104[5] , \R_DATA_TEMPR104[4] , 
        \R_DATA_TEMPR104[3] , \R_DATA_TEMPR104[2] , 
        \R_DATA_TEMPR104[1] , \R_DATA_TEMPR104[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[104][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[26] , \BLKY1[0] , \BLKY0[0] }), 
        .A_CLK(CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], 
        W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], 
        W_DATA[31], W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], 
        W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], 
        W_DATA[21], W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], 
        WBYTE_EN[2]}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], 
        W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], 
        W_ADDR[0], GND, GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[26] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA[19], 
        W_DATA[18], W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], 
        W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], W_DATA[9], 
        W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], 
        W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1126 (.A(\R_DATA_TEMPR60[33] ), .B(\R_DATA_TEMPR61[33] ), 
        .C(\R_DATA_TEMPR62[33] ), .D(\R_DATA_TEMPR63[33] ), .Y(
        OR4_1126_Y));
    OR4 OR4_951 (.A(\R_DATA_TEMPR24[29] ), .B(\R_DATA_TEMPR25[29] ), 
        .C(\R_DATA_TEMPR26[29] ), .D(\R_DATA_TEMPR27[29] ), .Y(
        OR4_951_Y));
    OR4 OR4_1510 (.A(\R_DATA_TEMPR12[3] ), .B(\R_DATA_TEMPR13[3] ), .C(
        \R_DATA_TEMPR14[3] ), .D(\R_DATA_TEMPR15[3] ), .Y(OR4_1510_Y));
    OR4 OR4_1465 (.A(\R_DATA_TEMPR20[29] ), .B(\R_DATA_TEMPR21[29] ), 
        .C(\R_DATA_TEMPR22[29] ), .D(\R_DATA_TEMPR23[29] ), .Y(
        OR4_1465_Y));
    OR4 OR4_1421 (.A(OR4_4_Y), .B(OR4_591_Y), .C(OR4_1384_Y), .D(
        OR4_1635_Y), .Y(OR4_1421_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[28]  (.A(CFG3_18_Y), .B(
        CFG3_3_Y), .Y(\BLKY2[28] ));
    OR4 OR4_642 (.A(\R_DATA_TEMPR92[4] ), .B(\R_DATA_TEMPR93[4] ), .C(
        \R_DATA_TEMPR94[4] ), .D(\R_DATA_TEMPR95[4] ), .Y(OR4_642_Y));
    OR4 OR4_1294 (.A(\R_DATA_TEMPR108[21] ), .B(\R_DATA_TEMPR109[21] ), 
        .C(\R_DATA_TEMPR110[21] ), .D(\R_DATA_TEMPR111[21] ), .Y(
        OR4_1294_Y));
    OR4 OR4_1509 (.A(OR4_1272_Y), .B(OR4_1132_Y), .C(OR4_1112_Y), .D(
        OR4_796_Y), .Y(OR4_1509_Y));
    OR2 OR2_30 (.A(\R_DATA_TEMPR84[20] ), .B(\R_DATA_TEMPR85[20] ), .Y(
        OR2_30_Y));
    OR4 OR4_1221 (.A(OR4_210_Y), .B(OR4_1418_Y), .C(OR4_1388_Y), .D(
        OR4_536_Y), .Y(OR4_1221_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%65%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R65C0 (.A_DOUT({
        \R_DATA_TEMPR65[39] , \R_DATA_TEMPR65[38] , 
        \R_DATA_TEMPR65[37] , \R_DATA_TEMPR65[36] , 
        \R_DATA_TEMPR65[35] , \R_DATA_TEMPR65[34] , 
        \R_DATA_TEMPR65[33] , \R_DATA_TEMPR65[32] , 
        \R_DATA_TEMPR65[31] , \R_DATA_TEMPR65[30] , 
        \R_DATA_TEMPR65[29] , \R_DATA_TEMPR65[28] , 
        \R_DATA_TEMPR65[27] , \R_DATA_TEMPR65[26] , 
        \R_DATA_TEMPR65[25] , \R_DATA_TEMPR65[24] , 
        \R_DATA_TEMPR65[23] , \R_DATA_TEMPR65[22] , 
        \R_DATA_TEMPR65[21] , \R_DATA_TEMPR65[20] }), .B_DOUT({
        \R_DATA_TEMPR65[19] , \R_DATA_TEMPR65[18] , 
        \R_DATA_TEMPR65[17] , \R_DATA_TEMPR65[16] , 
        \R_DATA_TEMPR65[15] , \R_DATA_TEMPR65[14] , 
        \R_DATA_TEMPR65[13] , \R_DATA_TEMPR65[12] , 
        \R_DATA_TEMPR65[11] , \R_DATA_TEMPR65[10] , 
        \R_DATA_TEMPR65[9] , \R_DATA_TEMPR65[8] , \R_DATA_TEMPR65[7] , 
        \R_DATA_TEMPR65[6] , \R_DATA_TEMPR65[5] , \R_DATA_TEMPR65[4] , 
        \R_DATA_TEMPR65[3] , \R_DATA_TEMPR65[2] , \R_DATA_TEMPR65[1] , 
        \R_DATA_TEMPR65[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[65][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[16] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[16] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_324 (.A(OR4_1334_Y), .B(OR4_829_Y), .C(OR4_888_Y), .D(
        OR4_1534_Y), .Y(OR4_324_Y));
    OR4 OR4_265 (.A(OR4_1091_Y), .B(OR4_834_Y), .C(OR4_559_Y), .D(
        OR4_1504_Y), .Y(OR4_265_Y));
    OR4 OR4_1397 (.A(\R_DATA_TEMPR0[2] ), .B(\R_DATA_TEMPR1[2] ), .C(
        \R_DATA_TEMPR2[2] ), .D(\R_DATA_TEMPR3[2] ), .Y(OR4_1397_Y));
    OR4 OR4_1128 (.A(OR4_446_Y), .B(OR4_127_Y), .C(OR4_110_Y), .D(
        OR4_897_Y), .Y(OR4_1128_Y));
    OR4 OR4_49 (.A(\R_DATA_TEMPR112[38] ), .B(\R_DATA_TEMPR113[38] ), 
        .C(\R_DATA_TEMPR114[38] ), .D(\R_DATA_TEMPR115[38] ), .Y(
        OR4_49_Y));
    OR4 OR4_599 (.A(\R_DATA_TEMPR0[23] ), .B(\R_DATA_TEMPR1[23] ), .C(
        \R_DATA_TEMPR2[23] ), .D(\R_DATA_TEMPR3[23] ), .Y(OR4_599_Y));
    OR2 OR2_14 (.A(\R_DATA_TEMPR84[14] ), .B(\R_DATA_TEMPR85[14] ), .Y(
        OR2_14_Y));
    OR2 OR2_37 (.A(\R_DATA_TEMPR84[12] ), .B(\R_DATA_TEMPR85[12] ), .Y(
        OR2_37_Y));
    OR4 OR4_1218 (.A(\R_DATA_TEMPR96[28] ), .B(\R_DATA_TEMPR97[28] ), 
        .C(\R_DATA_TEMPR98[28] ), .D(\R_DATA_TEMPR99[28] ), .Y(
        OR4_1218_Y));
    OR4 OR4_862 (.A(\R_DATA_TEMPR76[37] ), .B(\R_DATA_TEMPR77[37] ), 
        .C(\R_DATA_TEMPR78[37] ), .D(\R_DATA_TEMPR79[37] ), .Y(
        OR4_862_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%99%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R99C0 (.A_DOUT({
        \R_DATA_TEMPR99[39] , \R_DATA_TEMPR99[38] , 
        \R_DATA_TEMPR99[37] , \R_DATA_TEMPR99[36] , 
        \R_DATA_TEMPR99[35] , \R_DATA_TEMPR99[34] , 
        \R_DATA_TEMPR99[33] , \R_DATA_TEMPR99[32] , 
        \R_DATA_TEMPR99[31] , \R_DATA_TEMPR99[30] , 
        \R_DATA_TEMPR99[29] , \R_DATA_TEMPR99[28] , 
        \R_DATA_TEMPR99[27] , \R_DATA_TEMPR99[26] , 
        \R_DATA_TEMPR99[25] , \R_DATA_TEMPR99[24] , 
        \R_DATA_TEMPR99[23] , \R_DATA_TEMPR99[22] , 
        \R_DATA_TEMPR99[21] , \R_DATA_TEMPR99[20] }), .B_DOUT({
        \R_DATA_TEMPR99[19] , \R_DATA_TEMPR99[18] , 
        \R_DATA_TEMPR99[17] , \R_DATA_TEMPR99[16] , 
        \R_DATA_TEMPR99[15] , \R_DATA_TEMPR99[14] , 
        \R_DATA_TEMPR99[13] , \R_DATA_TEMPR99[12] , 
        \R_DATA_TEMPR99[11] , \R_DATA_TEMPR99[10] , 
        \R_DATA_TEMPR99[9] , \R_DATA_TEMPR99[8] , \R_DATA_TEMPR99[7] , 
        \R_DATA_TEMPR99[6] , \R_DATA_TEMPR99[5] , \R_DATA_TEMPR99[4] , 
        \R_DATA_TEMPR99[3] , \R_DATA_TEMPR99[2] , \R_DATA_TEMPR99[1] , 
        \R_DATA_TEMPR99[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[99][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[24] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[24] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%21%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C0 (.A_DOUT({
        \R_DATA_TEMPR21[39] , \R_DATA_TEMPR21[38] , 
        \R_DATA_TEMPR21[37] , \R_DATA_TEMPR21[36] , 
        \R_DATA_TEMPR21[35] , \R_DATA_TEMPR21[34] , 
        \R_DATA_TEMPR21[33] , \R_DATA_TEMPR21[32] , 
        \R_DATA_TEMPR21[31] , \R_DATA_TEMPR21[30] , 
        \R_DATA_TEMPR21[29] , \R_DATA_TEMPR21[28] , 
        \R_DATA_TEMPR21[27] , \R_DATA_TEMPR21[26] , 
        \R_DATA_TEMPR21[25] , \R_DATA_TEMPR21[24] , 
        \R_DATA_TEMPR21[23] , \R_DATA_TEMPR21[22] , 
        \R_DATA_TEMPR21[21] , \R_DATA_TEMPR21[20] }), .B_DOUT({
        \R_DATA_TEMPR21[19] , \R_DATA_TEMPR21[18] , 
        \R_DATA_TEMPR21[17] , \R_DATA_TEMPR21[16] , 
        \R_DATA_TEMPR21[15] , \R_DATA_TEMPR21[14] , 
        \R_DATA_TEMPR21[13] , \R_DATA_TEMPR21[12] , 
        \R_DATA_TEMPR21[11] , \R_DATA_TEMPR21[10] , 
        \R_DATA_TEMPR21[9] , \R_DATA_TEMPR21[8] , \R_DATA_TEMPR21[7] , 
        \R_DATA_TEMPR21[6] , \R_DATA_TEMPR21[5] , \R_DATA_TEMPR21[4] , 
        \R_DATA_TEMPR21[3] , \R_DATA_TEMPR21[2] , \R_DATA_TEMPR21[1] , 
        \R_DATA_TEMPR21[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[23]  (.A(CFG3_21_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[23] ));
    OR4 OR4_590 (.A(\R_DATA_TEMPR96[30] ), .B(\R_DATA_TEMPR97[30] ), 
        .C(\R_DATA_TEMPR98[30] ), .D(\R_DATA_TEMPR99[30] ), .Y(
        OR4_590_Y));
    OR4 OR4_121 (.A(\R_DATA_TEMPR20[32] ), .B(\R_DATA_TEMPR21[32] ), 
        .C(\R_DATA_TEMPR22[32] ), .D(\R_DATA_TEMPR23[32] ), .Y(
        OR4_121_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[5]  (.A(CFG3_22_Y), .B(
        CFG3_12_Y), .Y(\BLKX2[5] ));
    OR4 OR4_1183 (.A(\R_DATA_TEMPR52[4] ), .B(\R_DATA_TEMPR53[4] ), .C(
        \R_DATA_TEMPR54[4] ), .D(\R_DATA_TEMPR55[4] ), .Y(OR4_1183_Y));
    OR4 OR4_1142 (.A(OR4_998_Y), .B(OR4_405_Y), .C(OR4_644_Y), .D(
        OR4_1222_Y), .Y(OR4_1142_Y));
    OR4 OR4_919 (.A(\R_DATA_TEMPR40[22] ), .B(\R_DATA_TEMPR41[22] ), 
        .C(\R_DATA_TEMPR42[22] ), .D(\R_DATA_TEMPR43[22] ), .Y(
        OR4_919_Y));
    OR4 OR4_910 (.A(\R_DATA_TEMPR68[12] ), .B(\R_DATA_TEMPR69[12] ), 
        .C(\R_DATA_TEMPR70[12] ), .D(\R_DATA_TEMPR71[12] ), .Y(
        OR4_910_Y));
    OR4 \OR4_R_DATA[18]  (.A(OR4_1554_Y), .B(OR4_1343_Y), .C(OR4_597_Y)
        , .D(OR4_816_Y), .Y(R_DATA[18]));
    OR4 OR4_830 (.A(\R_DATA_TEMPR56[3] ), .B(\R_DATA_TEMPR57[3] ), .C(
        \R_DATA_TEMPR58[3] ), .D(\R_DATA_TEMPR59[3] ), .Y(OR4_830_Y));
    OR4 OR4_1177 (.A(\R_DATA_TEMPR72[8] ), .B(\R_DATA_TEMPR73[8] ), .C(
        \R_DATA_TEMPR74[8] ), .D(\R_DATA_TEMPR75[8] ), .Y(OR4_1177_Y));
    OR4 OR4_680 (.A(\R_DATA_TEMPR48[13] ), .B(\R_DATA_TEMPR49[13] ), 
        .C(\R_DATA_TEMPR50[13] ), .D(\R_DATA_TEMPR51[13] ), .Y(
        OR4_680_Y));
    OR4 OR4_113 (.A(OR4_1019_Y), .B(OR4_857_Y), .C(OR4_255_Y), .D(
        OR4_774_Y), .Y(OR4_113_Y));
    OR4 OR4_132 (.A(\R_DATA_TEMPR32[16] ), .B(\R_DATA_TEMPR33[16] ), 
        .C(\R_DATA_TEMPR34[16] ), .D(\R_DATA_TEMPR35[16] ), .Y(
        OR4_132_Y));
    OR4 OR4_7 (.A(\R_DATA_TEMPR96[36] ), .B(\R_DATA_TEMPR97[36] ), .C(
        \R_DATA_TEMPR98[36] ), .D(\R_DATA_TEMPR99[36] ), .Y(OR4_7_Y));
    OR4 OR4_1589 (.A(\R_DATA_TEMPR32[28] ), .B(\R_DATA_TEMPR33[28] ), 
        .C(\R_DATA_TEMPR34[28] ), .D(\R_DATA_TEMPR35[28] ), .Y(
        OR4_1589_Y));
    OR4 OR4_845 (.A(\R_DATA_TEMPR4[17] ), .B(\R_DATA_TEMPR5[17] ), .C(
        \R_DATA_TEMPR6[17] ), .D(\R_DATA_TEMPR7[17] ), .Y(OR4_845_Y));
    OR4 OR4_421 (.A(\R_DATA_TEMPR92[23] ), .B(\R_DATA_TEMPR93[23] ), 
        .C(\R_DATA_TEMPR94[23] ), .D(\R_DATA_TEMPR95[23] ), .Y(
        OR4_421_Y));
    OR4 OR4_935 (.A(\R_DATA_TEMPR36[34] ), .B(\R_DATA_TEMPR37[34] ), 
        .C(\R_DATA_TEMPR38[34] ), .D(\R_DATA_TEMPR39[34] ), .Y(
        OR4_935_Y));
    OR4 OR4_463 (.A(\R_DATA_TEMPR28[21] ), .B(\R_DATA_TEMPR29[21] ), 
        .C(\R_DATA_TEMPR30[21] ), .D(\R_DATA_TEMPR31[21] ), .Y(
        OR4_463_Y));
    OR4 OR4_755 (.A(\R_DATA_TEMPR52[39] ), .B(\R_DATA_TEMPR53[39] ), 
        .C(\R_DATA_TEMPR54[39] ), .D(\R_DATA_TEMPR55[39] ), .Y(
        OR4_755_Y));
    OR4 OR4_661 (.A(\R_DATA_TEMPR96[23] ), .B(\R_DATA_TEMPR97[23] ), 
        .C(\R_DATA_TEMPR98[23] ), .D(\R_DATA_TEMPR99[23] ), .Y(
        OR4_661_Y));
    OR4 OR4_657 (.A(\R_DATA_TEMPR116[5] ), .B(\R_DATA_TEMPR117[5] ), 
        .C(\R_DATA_TEMPR118[5] ), .D(\R_DATA_TEMPR119[5] ), .Y(
        OR4_657_Y));
    OR4 OR4_428 (.A(OR4_1412_Y), .B(OR4_1223_Y), .C(OR4_621_Y), .D(
        OR4_1134_Y), .Y(OR4_428_Y));
    OR4 OR4_1366 (.A(\R_DATA_TEMPR88[20] ), .B(\R_DATA_TEMPR89[20] ), 
        .C(\R_DATA_TEMPR90[20] ), .D(\R_DATA_TEMPR91[20] ), .Y(
        OR4_1366_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%103%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R103C0 (.A_DOUT({
        \R_DATA_TEMPR103[39] , \R_DATA_TEMPR103[38] , 
        \R_DATA_TEMPR103[37] , \R_DATA_TEMPR103[36] , 
        \R_DATA_TEMPR103[35] , \R_DATA_TEMPR103[34] , 
        \R_DATA_TEMPR103[33] , \R_DATA_TEMPR103[32] , 
        \R_DATA_TEMPR103[31] , \R_DATA_TEMPR103[30] , 
        \R_DATA_TEMPR103[29] , \R_DATA_TEMPR103[28] , 
        \R_DATA_TEMPR103[27] , \R_DATA_TEMPR103[26] , 
        \R_DATA_TEMPR103[25] , \R_DATA_TEMPR103[24] , 
        \R_DATA_TEMPR103[23] , \R_DATA_TEMPR103[22] , 
        \R_DATA_TEMPR103[21] , \R_DATA_TEMPR103[20] }), .B_DOUT({
        \R_DATA_TEMPR103[19] , \R_DATA_TEMPR103[18] , 
        \R_DATA_TEMPR103[17] , \R_DATA_TEMPR103[16] , 
        \R_DATA_TEMPR103[15] , \R_DATA_TEMPR103[14] , 
        \R_DATA_TEMPR103[13] , \R_DATA_TEMPR103[12] , 
        \R_DATA_TEMPR103[11] , \R_DATA_TEMPR103[10] , 
        \R_DATA_TEMPR103[9] , \R_DATA_TEMPR103[8] , 
        \R_DATA_TEMPR103[7] , \R_DATA_TEMPR103[6] , 
        \R_DATA_TEMPR103[5] , \R_DATA_TEMPR103[4] , 
        \R_DATA_TEMPR103[3] , \R_DATA_TEMPR103[2] , 
        \R_DATA_TEMPR103[1] , \R_DATA_TEMPR103[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[103][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[25] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[25] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1453 (.A(\R_DATA_TEMPR60[12] ), .B(\R_DATA_TEMPR61[12] ), 
        .C(\R_DATA_TEMPR62[12] ), .D(\R_DATA_TEMPR63[12] ), .Y(
        OR4_1453_Y));
    OR4 OR4_756 (.A(\R_DATA_TEMPR4[28] ), .B(\R_DATA_TEMPR5[28] ), .C(
        \R_DATA_TEMPR6[28] ), .D(\R_DATA_TEMPR7[28] ), .Y(OR4_756_Y));
    OR4 OR4_268 (.A(\R_DATA_TEMPR88[1] ), .B(\R_DATA_TEMPR89[1] ), .C(
        \R_DATA_TEMPR90[1] ), .D(\R_DATA_TEMPR91[1] ), .Y(OR4_268_Y));
    OR4 OR4_387 (.A(\R_DATA_TEMPR100[0] ), .B(\R_DATA_TEMPR101[0] ), 
        .C(\R_DATA_TEMPR102[0] ), .D(\R_DATA_TEMPR103[0] ), .Y(
        OR4_387_Y));
    OR4 OR4_180 (.A(\R_DATA_TEMPR96[29] ), .B(\R_DATA_TEMPR97[29] ), 
        .C(\R_DATA_TEMPR98[29] ), .D(\R_DATA_TEMPR99[29] ), .Y(
        OR4_180_Y));
    OR4 OR4_1495 (.A(\R_DATA_TEMPR48[2] ), .B(\R_DATA_TEMPR49[2] ), .C(
        \R_DATA_TEMPR50[2] ), .D(\R_DATA_TEMPR51[2] ), .Y(OR4_1495_Y));
    OR4 OR4_105 (.A(\R_DATA_TEMPR60[15] ), .B(\R_DATA_TEMPR61[15] ), 
        .C(\R_DATA_TEMPR62[15] ), .D(\R_DATA_TEMPR63[15] ), .Y(
        OR4_105_Y));
    OR4 OR4_788 (.A(\R_DATA_TEMPR52[16] ), .B(\R_DATA_TEMPR53[16] ), 
        .C(\R_DATA_TEMPR54[16] ), .D(\R_DATA_TEMPR55[16] ), .Y(
        OR4_788_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%95%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R95C0 (.A_DOUT({
        \R_DATA_TEMPR95[39] , \R_DATA_TEMPR95[38] , 
        \R_DATA_TEMPR95[37] , \R_DATA_TEMPR95[36] , 
        \R_DATA_TEMPR95[35] , \R_DATA_TEMPR95[34] , 
        \R_DATA_TEMPR95[33] , \R_DATA_TEMPR95[32] , 
        \R_DATA_TEMPR95[31] , \R_DATA_TEMPR95[30] , 
        \R_DATA_TEMPR95[29] , \R_DATA_TEMPR95[28] , 
        \R_DATA_TEMPR95[27] , \R_DATA_TEMPR95[26] , 
        \R_DATA_TEMPR95[25] , \R_DATA_TEMPR95[24] , 
        \R_DATA_TEMPR95[23] , \R_DATA_TEMPR95[22] , 
        \R_DATA_TEMPR95[21] , \R_DATA_TEMPR95[20] }), .B_DOUT({
        \R_DATA_TEMPR95[19] , \R_DATA_TEMPR95[18] , 
        \R_DATA_TEMPR95[17] , \R_DATA_TEMPR95[16] , 
        \R_DATA_TEMPR95[15] , \R_DATA_TEMPR95[14] , 
        \R_DATA_TEMPR95[13] , \R_DATA_TEMPR95[12] , 
        \R_DATA_TEMPR95[11] , \R_DATA_TEMPR95[10] , 
        \R_DATA_TEMPR95[9] , \R_DATA_TEMPR95[8] , \R_DATA_TEMPR95[7] , 
        \R_DATA_TEMPR95[6] , \R_DATA_TEMPR95[5] , \R_DATA_TEMPR95[4] , 
        \R_DATA_TEMPR95[3] , \R_DATA_TEMPR95[2] , \R_DATA_TEMPR95[1] , 
        \R_DATA_TEMPR95[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[95][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[23] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[23] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_407 (.A(\R_DATA_TEMPR4[8] ), .B(\R_DATA_TEMPR5[8] ), .C(
        \R_DATA_TEMPR6[8] ), .D(\R_DATA_TEMPR7[8] ), .Y(OR4_407_Y));
    OR4 OR4_1505 (.A(OR4_427_Y), .B(OR4_700_Y), .C(OR4_691_Y), .D(
        OR4_960_Y), .Y(OR4_1505_Y));
    CFG3 #( .INIT(8'h10) )  CFG3_15 (.A(R_ADDR[13]), .B(R_ADDR[12]), 
        .C(R_ADDR[11]), .Y(CFG3_15_Y));
    OR4 OR4_175 (.A(\R_DATA_TEMPR72[19] ), .B(\R_DATA_TEMPR73[19] ), 
        .C(\R_DATA_TEMPR74[19] ), .D(\R_DATA_TEMPR75[19] ), .Y(
        OR4_175_Y));
    OR4 OR4_393 (.A(\R_DATA_TEMPR36[22] ), .B(\R_DATA_TEMPR37[22] ), 
        .C(\R_DATA_TEMPR38[22] ), .D(\R_DATA_TEMPR39[22] ), .Y(
        OR4_393_Y));
    OR4 OR4_790 (.A(\R_DATA_TEMPR48[37] ), .B(\R_DATA_TEMPR49[37] ), 
        .C(\R_DATA_TEMPR50[37] ), .D(\R_DATA_TEMPR51[37] ), .Y(
        OR4_790_Y));
    OR4 OR4_1619 (.A(\R_DATA_TEMPR40[5] ), .B(\R_DATA_TEMPR41[5] ), .C(
        \R_DATA_TEMPR42[5] ), .D(\R_DATA_TEMPR43[5] ), .Y(OR4_1619_Y));
    OR4 OR4_1115 (.A(\R_DATA_TEMPR4[20] ), .B(\R_DATA_TEMPR5[20] ), .C(
        \R_DATA_TEMPR6[20] ), .D(\R_DATA_TEMPR7[20] ), .Y(OR4_1115_Y));
    OR4 OR4_239 (.A(\R_DATA_TEMPR28[28] ), .B(\R_DATA_TEMPR29[28] ), 
        .C(\R_DATA_TEMPR30[28] ), .D(\R_DATA_TEMPR31[28] ), .Y(
        OR4_239_Y));
    OR4 OR4_42 (.A(OR4_1225_Y), .B(OR4_1261_Y), .C(OR4_164_Y), .D(
        OR4_1191_Y), .Y(OR4_42_Y));
    OR4 OR4_529 (.A(OR4_852_Y), .B(OR4_264_Y), .C(OR4_789_Y), .D(
        OR4_1246_Y), .Y(OR4_529_Y));
    OR4 OR4_477 (.A(\R_DATA_TEMPR112[37] ), .B(\R_DATA_TEMPR113[37] ), 
        .C(\R_DATA_TEMPR114[37] ), .D(\R_DATA_TEMPR115[37] ), .Y(
        OR4_477_Y));
    OR4 OR4_1206 (.A(\R_DATA_TEMPR116[8] ), .B(\R_DATA_TEMPR117[8] ), 
        .C(\R_DATA_TEMPR118[8] ), .D(\R_DATA_TEMPR119[8] ), .Y(
        OR4_1206_Y));
    OR4 OR4_1011 (.A(OR4_458_Y), .B(OR4_279_Y), .C(OR4_1317_Y), .D(
        OR4_195_Y), .Y(OR4_1011_Y));
    OR4 OR4_492 (.A(\R_DATA_TEMPR88[18] ), .B(\R_DATA_TEMPR89[18] ), 
        .C(\R_DATA_TEMPR90[18] ), .D(\R_DATA_TEMPR91[18] ), .Y(
        OR4_492_Y));
    OR4 OR4_520 (.A(\R_DATA_TEMPR40[11] ), .B(\R_DATA_TEMPR41[11] ), 
        .C(\R_DATA_TEMPR42[11] ), .D(\R_DATA_TEMPR43[11] ), .Y(
        OR4_520_Y));
    OR4 OR4_499 (.A(OR4_1411_Y), .B(OR4_76_Y), .C(OR4_1145_Y), .D(
        OR4_379_Y), .Y(OR4_499_Y));
    OR4 OR4_88 (.A(\R_DATA_TEMPR64[17] ), .B(\R_DATA_TEMPR65[17] ), .C(
        \R_DATA_TEMPR66[17] ), .D(\R_DATA_TEMPR67[17] ), .Y(OR4_88_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[7]  (.A(CFG3_23_Y), .B(
        CFG3_12_Y), .Y(\BLKX2[7] ));
    OR4 OR4_1308 (.A(\R_DATA_TEMPR24[17] ), .B(\R_DATA_TEMPR25[17] ), 
        .C(\R_DATA_TEMPR26[17] ), .D(\R_DATA_TEMPR27[17] ), .Y(
        OR4_1308_Y));
    OR4 OR4_205 (.A(\R_DATA_TEMPR28[35] ), .B(\R_DATA_TEMPR29[35] ), 
        .C(\R_DATA_TEMPR30[35] ), .D(\R_DATA_TEMPR31[35] ), .Y(
        OR4_205_Y));
    OR4 OR4_887 (.A(\R_DATA_TEMPR100[9] ), .B(\R_DATA_TEMPR101[9] ), 
        .C(\R_DATA_TEMPR102[9] ), .D(\R_DATA_TEMPR103[9] ), .Y(
        OR4_887_Y));
    OR4 OR4_188 (.A(OR4_256_Y), .B(OR4_372_Y), .C(OR4_357_Y), .D(
        OR4_18_Y), .Y(OR4_188_Y));
    OR4 OR4_984 (.A(\R_DATA_TEMPR108[20] ), .B(\R_DATA_TEMPR109[20] ), 
        .C(\R_DATA_TEMPR110[20] ), .D(\R_DATA_TEMPR111[20] ), .Y(
        OR4_984_Y));
    OR4 OR4_810 (.A(\R_DATA_TEMPR32[25] ), .B(\R_DATA_TEMPR33[25] ), 
        .C(\R_DATA_TEMPR34[25] ), .D(\R_DATA_TEMPR35[25] ), .Y(
        OR4_810_Y));
    OR4 OR4_196 (.A(OR4_574_Y), .B(OR4_1136_Y), .C(OR4_317_Y), .D(
        OR4_565_Y), .Y(OR4_196_Y));
    OR4 OR4_802 (.A(\R_DATA_TEMPR24[26] ), .B(\R_DATA_TEMPR25[26] ), 
        .C(\R_DATA_TEMPR26[26] ), .D(\R_DATA_TEMPR27[26] ), .Y(
        OR4_802_Y));
    OR4 OR4_1468 (.A(\R_DATA_TEMPR8[33] ), .B(\R_DATA_TEMPR9[33] ), .C(
        \R_DATA_TEMPR10[33] ), .D(\R_DATA_TEMPR11[33] ), .Y(OR4_1468_Y)
        );
    OR4 OR4_112 (.A(\R_DATA_TEMPR104[31] ), .B(\R_DATA_TEMPR105[31] ), 
        .C(\R_DATA_TEMPR106[31] ), .D(\R_DATA_TEMPR107[31] ), .Y(
        OR4_112_Y));
    OR4 OR4_275 (.A(OR4_745_Y), .B(OR4_491_Y), .C(OR4_201_Y), .D(
        OR4_570_Y), .Y(OR4_275_Y));
    OR4 OR4_1633 (.A(\R_DATA_TEMPR44[8] ), .B(\R_DATA_TEMPR45[8] ), .C(
        \R_DATA_TEMPR46[8] ), .D(\R_DATA_TEMPR47[8] ), .Y(OR4_1633_Y));
    OR4 OR4_1270 (.A(\R_DATA_TEMPR44[30] ), .B(\R_DATA_TEMPR45[30] ), 
        .C(\R_DATA_TEMPR46[30] ), .D(\R_DATA_TEMPR47[30] ), .Y(
        OR4_1270_Y));
    OR4 OR4_1013 (.A(\R_DATA_TEMPR4[35] ), .B(\R_DATA_TEMPR5[35] ), .C(
        \R_DATA_TEMPR6[35] ), .D(\R_DATA_TEMPR7[35] ), .Y(OR4_1013_Y));
    OR4 OR4_915 (.A(\R_DATA_TEMPR4[1] ), .B(\R_DATA_TEMPR5[1] ), .C(
        \R_DATA_TEMPR6[1] ), .D(\R_DATA_TEMPR7[1] ), .Y(OR4_915_Y));
    OR4 OR4_839 (.A(\R_DATA_TEMPR60[16] ), .B(\R_DATA_TEMPR61[16] ), 
        .C(\R_DATA_TEMPR62[16] ), .D(\R_DATA_TEMPR63[16] ), .Y(
        OR4_839_Y));
    OR4 OR4_1585 (.A(\R_DATA_TEMPR0[8] ), .B(\R_DATA_TEMPR1[8] ), .C(
        \R_DATA_TEMPR2[8] ), .D(\R_DATA_TEMPR3[8] ), .Y(OR4_1585_Y));
    OR4 OR4_1396 (.A(\R_DATA_TEMPR52[3] ), .B(\R_DATA_TEMPR53[3] ), .C(
        \R_DATA_TEMPR54[3] ), .D(\R_DATA_TEMPR55[3] ), .Y(OR4_1396_Y));
    OR4 OR4_872 (.A(\R_DATA_TEMPR104[36] ), .B(\R_DATA_TEMPR105[36] ), 
        .C(\R_DATA_TEMPR106[36] ), .D(\R_DATA_TEMPR107[36] ), .Y(
        OR4_872_Y));
    OR4 OR4_646 (.A(OR4_1385_Y), .B(OR4_56_Y), .C(OR4_307_Y), .D(
        OR4_105_Y), .Y(OR4_646_Y));
    OR4 OR4_1412 (.A(\R_DATA_TEMPR96[39] ), .B(\R_DATA_TEMPR97[39] ), 
        .C(\R_DATA_TEMPR98[39] ), .D(\R_DATA_TEMPR99[39] ), .Y(
        OR4_1412_Y));
    OR4 \OR4_R_DATA[37]  (.A(OR4_724_Y), .B(OR4_1509_Y), .C(OR4_297_Y), 
        .D(OR4_445_Y), .Y(R_DATA[37]));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%116%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R116C0 (.A_DOUT({
        \R_DATA_TEMPR116[39] , \R_DATA_TEMPR116[38] , 
        \R_DATA_TEMPR116[37] , \R_DATA_TEMPR116[36] , 
        \R_DATA_TEMPR116[35] , \R_DATA_TEMPR116[34] , 
        \R_DATA_TEMPR116[33] , \R_DATA_TEMPR116[32] , 
        \R_DATA_TEMPR116[31] , \R_DATA_TEMPR116[30] , 
        \R_DATA_TEMPR116[29] , \R_DATA_TEMPR116[28] , 
        \R_DATA_TEMPR116[27] , \R_DATA_TEMPR116[26] , 
        \R_DATA_TEMPR116[25] , \R_DATA_TEMPR116[24] , 
        \R_DATA_TEMPR116[23] , \R_DATA_TEMPR116[22] , 
        \R_DATA_TEMPR116[21] , \R_DATA_TEMPR116[20] }), .B_DOUT({
        \R_DATA_TEMPR116[19] , \R_DATA_TEMPR116[18] , 
        \R_DATA_TEMPR116[17] , \R_DATA_TEMPR116[16] , 
        \R_DATA_TEMPR116[15] , \R_DATA_TEMPR116[14] , 
        \R_DATA_TEMPR116[13] , \R_DATA_TEMPR116[12] , 
        \R_DATA_TEMPR116[11] , \R_DATA_TEMPR116[10] , 
        \R_DATA_TEMPR116[9] , \R_DATA_TEMPR116[8] , 
        \R_DATA_TEMPR116[7] , \R_DATA_TEMPR116[6] , 
        \R_DATA_TEMPR116[5] , \R_DATA_TEMPR116[4] , 
        \R_DATA_TEMPR116[3] , \R_DATA_TEMPR116[2] , 
        \R_DATA_TEMPR116[1] , \R_DATA_TEMPR116[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[116][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[29] , \BLKY1[0] , \BLKY0[0] }), 
        .A_CLK(CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], 
        W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], 
        W_DATA[31], W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], 
        W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], 
        W_DATA[21], W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], 
        WBYTE_EN[2]}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], 
        W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], 
        W_ADDR[0], GND, GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[29] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA[19], 
        W_DATA[18], W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], 
        W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], W_DATA[9], 
        W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], 
        W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1534 (.A(\R_DATA_TEMPR76[35] ), .B(\R_DATA_TEMPR77[35] ), 
        .C(\R_DATA_TEMPR78[35] ), .D(\R_DATA_TEMPR79[35] ), .Y(
        OR4_1534_Y));
    OR4 OR4_1577 (.A(\R_DATA_TEMPR60[8] ), .B(\R_DATA_TEMPR61[8] ), .C(
        \R_DATA_TEMPR62[8] ), .D(\R_DATA_TEMPR63[8] ), .Y(OR4_1577_Y));
    OR4 OR4_1286 (.A(\R_DATA_TEMPR20[4] ), .B(\R_DATA_TEMPR21[4] ), .C(
        \R_DATA_TEMPR22[4] ), .D(\R_DATA_TEMPR23[4] ), .Y(OR4_1286_Y));
    OR4 OR4_257 (.A(\R_DATA_TEMPR32[33] ), .B(\R_DATA_TEMPR33[33] ), 
        .C(\R_DATA_TEMPR34[33] ), .D(\R_DATA_TEMPR35[33] ), .Y(
        OR4_257_Y));
    OR4 OR4_1372 (.A(\R_DATA_TEMPR104[4] ), .B(\R_DATA_TEMPR105[4] ), 
        .C(\R_DATA_TEMPR106[4] ), .D(\R_DATA_TEMPR107[4] ), .Y(
        OR4_1372_Y));
    OR4 OR4_398 (.A(OR4_496_Y), .B(OR4_1018_Y), .C(OR4_1450_Y), .D(
        OR4_553_Y), .Y(OR4_398_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%100%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R100C0 (.A_DOUT({
        \R_DATA_TEMPR100[39] , \R_DATA_TEMPR100[38] , 
        \R_DATA_TEMPR100[37] , \R_DATA_TEMPR100[36] , 
        \R_DATA_TEMPR100[35] , \R_DATA_TEMPR100[34] , 
        \R_DATA_TEMPR100[33] , \R_DATA_TEMPR100[32] , 
        \R_DATA_TEMPR100[31] , \R_DATA_TEMPR100[30] , 
        \R_DATA_TEMPR100[29] , \R_DATA_TEMPR100[28] , 
        \R_DATA_TEMPR100[27] , \R_DATA_TEMPR100[26] , 
        \R_DATA_TEMPR100[25] , \R_DATA_TEMPR100[24] , 
        \R_DATA_TEMPR100[23] , \R_DATA_TEMPR100[22] , 
        \R_DATA_TEMPR100[21] , \R_DATA_TEMPR100[20] }), .B_DOUT({
        \R_DATA_TEMPR100[19] , \R_DATA_TEMPR100[18] , 
        \R_DATA_TEMPR100[17] , \R_DATA_TEMPR100[16] , 
        \R_DATA_TEMPR100[15] , \R_DATA_TEMPR100[14] , 
        \R_DATA_TEMPR100[13] , \R_DATA_TEMPR100[12] , 
        \R_DATA_TEMPR100[11] , \R_DATA_TEMPR100[10] , 
        \R_DATA_TEMPR100[9] , \R_DATA_TEMPR100[8] , 
        \R_DATA_TEMPR100[7] , \R_DATA_TEMPR100[6] , 
        \R_DATA_TEMPR100[5] , \R_DATA_TEMPR100[4] , 
        \R_DATA_TEMPR100[3] , \R_DATA_TEMPR100[2] , 
        \R_DATA_TEMPR100[1] , \R_DATA_TEMPR100[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[100][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[25] , \BLKY1[0] , \BLKY0[0] }), 
        .A_CLK(CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], 
        W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], 
        W_DATA[31], W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], 
        W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], 
        W_DATA[21], W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], 
        WBYTE_EN[2]}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], 
        W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], 
        W_ADDR[0], GND, GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[25] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA[19], 
        W_DATA[18], W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], 
        W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], W_DATA[9], 
        W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], 
        W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1009 (.A(\R_DATA_TEMPR88[23] ), .B(\R_DATA_TEMPR89[23] ), 
        .C(\R_DATA_TEMPR90[23] ), .D(\R_DATA_TEMPR91[23] ), .Y(
        OR4_1009_Y));
    OR4 OR4_157 (.A(OR4_875_Y), .B(OR4_1106_Y), .C(OR4_1081_Y), .D(
        OR4_230_Y), .Y(OR4_157_Y));
    OR4 OR4_1335 (.A(\R_DATA_TEMPR76[15] ), .B(\R_DATA_TEMPR77[15] ), 
        .C(\R_DATA_TEMPR78[15] ), .D(\R_DATA_TEMPR79[15] ), .Y(
        OR4_1335_Y));
    OR4 OR4_1272 (.A(OR4_41_Y), .B(OR4_1165_Y), .C(OR4_1227_Y), .D(
        OR4_862_Y), .Y(OR4_1272_Y));
    OR4 OR4_561 (.A(OR4_662_Y), .B(OR4_935_Y), .C(OR4_916_Y), .D(
        OR4_604_Y), .Y(OR4_561_Y));
    OR4 OR4_403 (.A(OR4_475_Y), .B(OR4_325_Y), .C(OR4_442_Y), .D(
        OR4_976_Y), .Y(OR4_403_Y));
    OR4 OR4_1388 (.A(\R_DATA_TEMPR40[10] ), .B(\R_DATA_TEMPR41[10] ), 
        .C(\R_DATA_TEMPR42[10] ), .D(\R_DATA_TEMPR43[10] ), .Y(
        OR4_1388_Y));
    OR4 OR4_1153 (.A(\R_DATA_TEMPR80[36] ), .B(\R_DATA_TEMPR81[36] ), 
        .C(\R_DATA_TEMPR82[36] ), .D(\R_DATA_TEMPR83[36] ), .Y(
        OR4_1153_Y));
    OR4 OR4_601 (.A(\R_DATA_TEMPR56[25] ), .B(\R_DATA_TEMPR57[25] ), 
        .C(\R_DATA_TEMPR58[25] ), .D(\R_DATA_TEMPR59[25] ), .Y(
        OR4_601_Y));
    CFG3 #( .INIT(8'h80) )  CFG3_7 (.A(W_EN), .B(W_ADDR[15]), .C(
        W_ADDR[14]), .Y(CFG3_7_Y));
    OR4 OR4_1164 (.A(\R_DATA_TEMPR64[7] ), .B(\R_DATA_TEMPR65[7] ), .C(
        \R_DATA_TEMPR66[7] ), .D(\R_DATA_TEMPR67[7] ), .Y(OR4_1164_Y));
    OR4 OR4_208 (.A(\R_DATA_TEMPR24[30] ), .B(\R_DATA_TEMPR25[30] ), 
        .C(\R_DATA_TEMPR26[30] ), .D(\R_DATA_TEMPR27[30] ), .Y(
        OR4_208_Y));
    OR4 OR4_219 (.A(OR4_521_Y), .B(OR4_1448_Y), .C(OR4_908_Y), .D(
        OR4_365_Y), .Y(OR4_219_Y));
    OR4 \OR4_R_DATA[19]  (.A(OR4_527_Y), .B(OR4_157_Y), .C(OR4_47_Y), 
        .D(OR4_1415_Y), .Y(R_DATA[19]));
    OR4 OR4_323 (.A(OR4_930_Y), .B(OR4_1249_Y), .C(OR4_1496_Y), .D(
        OR4_1302_Y), .Y(OR4_323_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[19]  (.A(CFG3_19_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[19] ));
    OR4 OR4_720 (.A(\R_DATA_TEMPR12[36] ), .B(\R_DATA_TEMPR13[36] ), 
        .C(\R_DATA_TEMPR14[36] ), .D(\R_DATA_TEMPR15[36] ), .Y(
        OR4_720_Y));
    OR4 OR4_473 (.A(\R_DATA_TEMPR44[1] ), .B(\R_DATA_TEMPR45[1] ), .C(
        \R_DATA_TEMPR46[1] ), .D(\R_DATA_TEMPR47[1] ), .Y(OR4_473_Y));
    OR4 OR4_1474 (.A(OR4_90_Y), .B(OR2_26_Y), .C(\R_DATA_TEMPR86[27] ), 
        .D(\R_DATA_TEMPR87[27] ), .Y(OR4_1474_Y));
    OR4 OR4_671 (.A(\R_DATA_TEMPR8[4] ), .B(\R_DATA_TEMPR9[4] ), .C(
        \R_DATA_TEMPR10[4] ), .D(\R_DATA_TEMPR11[4] ), .Y(OR4_671_Y));
    OR4 OR4_1560 (.A(OR4_410_Y), .B(OR4_602_Y), .C(OR4_575_Y), .D(
        OR4_1356_Y), .Y(OR4_1560_Y));
    OR2 OR2_38 (.A(\R_DATA_TEMPR84[10] ), .B(\R_DATA_TEMPR85[10] ), .Y(
        OR2_38_Y));
    OR4 OR4_737 (.A(\R_DATA_TEMPR96[6] ), .B(\R_DATA_TEMPR97[6] ), .C(
        \R_DATA_TEMPR98[6] ), .D(\R_DATA_TEMPR99[6] ), .Y(OR4_737_Y));
    OR4 OR4_422 (.A(\R_DATA_TEMPR60[1] ), .B(\R_DATA_TEMPR61[1] ), .C(
        \R_DATA_TEMPR62[1] ), .D(\R_DATA_TEMPR63[1] ), .Y(OR4_422_Y));
    OR4 OR4_278 (.A(\R_DATA_TEMPR100[15] ), .B(\R_DATA_TEMPR101[15] ), 
        .C(\R_DATA_TEMPR102[15] ), .D(\R_DATA_TEMPR103[15] ), .Y(
        OR4_278_Y));
    OR4 OR4_1559 (.A(\R_DATA_TEMPR116[18] ), .B(\R_DATA_TEMPR117[18] ), 
        .C(\R_DATA_TEMPR118[18] ), .D(\R_DATA_TEMPR119[18] ), .Y(
        OR4_1559_Y));
    OR4 OR4_753 (.A(\R_DATA_TEMPR92[20] ), .B(\R_DATA_TEMPR93[20] ), 
        .C(\R_DATA_TEMPR94[20] ), .D(\R_DATA_TEMPR95[20] ), .Y(
        OR4_753_Y));
    OR4 OR4_734 (.A(\R_DATA_TEMPR24[15] ), .B(\R_DATA_TEMPR25[15] ), 
        .C(\R_DATA_TEMPR26[15] ), .D(\R_DATA_TEMPR27[15] ), .Y(
        OR4_734_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%72%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R72C0 (.A_DOUT({
        \R_DATA_TEMPR72[39] , \R_DATA_TEMPR72[38] , 
        \R_DATA_TEMPR72[37] , \R_DATA_TEMPR72[36] , 
        \R_DATA_TEMPR72[35] , \R_DATA_TEMPR72[34] , 
        \R_DATA_TEMPR72[33] , \R_DATA_TEMPR72[32] , 
        \R_DATA_TEMPR72[31] , \R_DATA_TEMPR72[30] , 
        \R_DATA_TEMPR72[29] , \R_DATA_TEMPR72[28] , 
        \R_DATA_TEMPR72[27] , \R_DATA_TEMPR72[26] , 
        \R_DATA_TEMPR72[25] , \R_DATA_TEMPR72[24] , 
        \R_DATA_TEMPR72[23] , \R_DATA_TEMPR72[22] , 
        \R_DATA_TEMPR72[21] , \R_DATA_TEMPR72[20] }), .B_DOUT({
        \R_DATA_TEMPR72[19] , \R_DATA_TEMPR72[18] , 
        \R_DATA_TEMPR72[17] , \R_DATA_TEMPR72[16] , 
        \R_DATA_TEMPR72[15] , \R_DATA_TEMPR72[14] , 
        \R_DATA_TEMPR72[13] , \R_DATA_TEMPR72[12] , 
        \R_DATA_TEMPR72[11] , \R_DATA_TEMPR72[10] , 
        \R_DATA_TEMPR72[9] , \R_DATA_TEMPR72[8] , \R_DATA_TEMPR72[7] , 
        \R_DATA_TEMPR72[6] , \R_DATA_TEMPR72[5] , \R_DATA_TEMPR72[4] , 
        \R_DATA_TEMPR72[3] , \R_DATA_TEMPR72[2] , \R_DATA_TEMPR72[1] , 
        \R_DATA_TEMPR72[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[72][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[18] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[18] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1274 (.A(\R_DATA_TEMPR12[33] ), .B(\R_DATA_TEMPR13[33] ), 
        .C(\R_DATA_TEMPR14[33] ), .D(\R_DATA_TEMPR15[33] ), .Y(
        OR4_1274_Y));
    OR4 OR4_1548 (.A(\R_DATA_TEMPR120[15] ), .B(\R_DATA_TEMPR121[15] ), 
        .C(\R_DATA_TEMPR122[15] ), .D(\R_DATA_TEMPR123[15] ), .Y(
        OR4_1548_Y));
    OR4 OR4_23 (.A(OR4_5_Y), .B(OR4_868_Y), .C(OR4_24_Y), .D(OR4_293_Y)
        , .Y(OR4_23_Y));
    OR4 OR4_199 (.A(\R_DATA_TEMPR12[6] ), .B(\R_DATA_TEMPR13[6] ), .C(
        \R_DATA_TEMPR14[6] ), .D(\R_DATA_TEMPR15[6] ), .Y(OR4_199_Y));
    OR4 OR4_254 (.A(\R_DATA_TEMPR28[7] ), .B(\R_DATA_TEMPR29[7] ), .C(
        \R_DATA_TEMPR30[7] ), .D(\R_DATA_TEMPR31[7] ), .Y(OR4_254_Y));
    OR4 OR4_1498 (.A(\R_DATA_TEMPR44[14] ), .B(\R_DATA_TEMPR45[14] ), 
        .C(\R_DATA_TEMPR46[14] ), .D(\R_DATA_TEMPR47[14] ), .Y(
        OR4_1498_Y));
    OR4 OR4_429 (.A(\R_DATA_TEMPR96[26] ), .B(\R_DATA_TEMPR97[26] ), 
        .C(\R_DATA_TEMPR98[26] ), .D(\R_DATA_TEMPR99[26] ), .Y(
        OR4_429_Y));
    OR4 OR4_1268 (.A(\R_DATA_TEMPR4[11] ), .B(\R_DATA_TEMPR5[11] ), .C(
        \R_DATA_TEMPR6[11] ), .D(\R_DATA_TEMPR7[11] ), .Y(OR4_1268_Y));
    OR4 OR4_262 (.A(\R_DATA_TEMPR100[32] ), .B(\R_DATA_TEMPR101[32] ), 
        .C(\R_DATA_TEMPR102[32] ), .D(\R_DATA_TEMPR103[32] ), .Y(
        OR4_262_Y));
    OR4 OR4_1377 (.A(\R_DATA_TEMPR8[8] ), .B(\R_DATA_TEMPR9[8] ), .C(
        \R_DATA_TEMPR10[8] ), .D(\R_DATA_TEMPR11[8] ), .Y(OR4_1377_Y));
    OR4 OR4_1249 (.A(\R_DATA_TEMPR100[16] ), .B(\R_DATA_TEMPR101[16] ), 
        .C(\R_DATA_TEMPR102[16] ), .D(\R_DATA_TEMPR103[16] ), .Y(
        OR4_1249_Y));
    OR4 OR4_1089 (.A(OR4_1258_Y), .B(OR4_1519_Y), .C(OR4_74_Y), .D(
        OR4_1275_Y), .Y(OR4_1089_Y));
    OR4 OR4_831 (.A(\R_DATA_TEMPR48[31] ), .B(\R_DATA_TEMPR49[31] ), 
        .C(\R_DATA_TEMPR50[31] ), .D(\R_DATA_TEMPR51[31] ), .Y(
        OR4_831_Y));
    OR4 OR4_126 (.A(\R_DATA_TEMPR88[33] ), .B(\R_DATA_TEMPR89[33] ), 
        .C(\R_DATA_TEMPR90[33] ), .D(\R_DATA_TEMPR91[33] ), .Y(
        OR4_126_Y));
    OR4 OR4_1623 (.A(\R_DATA_TEMPR4[25] ), .B(\R_DATA_TEMPR5[25] ), .C(
        \R_DATA_TEMPR6[25] ), .D(\R_DATA_TEMPR7[25] ), .Y(OR4_1623_Y));
    OR4 OR4_819 (.A(\R_DATA_TEMPR32[32] ), .B(\R_DATA_TEMPR33[32] ), 
        .C(\R_DATA_TEMPR34[32] ), .D(\R_DATA_TEMPR35[32] ), .Y(
        OR4_819_Y));
    OR4 OR4_94 (.A(\R_DATA_TEMPR124[17] ), .B(\R_DATA_TEMPR125[17] ), 
        .C(\R_DATA_TEMPR126[17] ), .D(\R_DATA_TEMPR127[17] ), .Y(
        OR4_94_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%82%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R82C0 (.A_DOUT({
        \R_DATA_TEMPR82[39] , \R_DATA_TEMPR82[38] , 
        \R_DATA_TEMPR82[37] , \R_DATA_TEMPR82[36] , 
        \R_DATA_TEMPR82[35] , \R_DATA_TEMPR82[34] , 
        \R_DATA_TEMPR82[33] , \R_DATA_TEMPR82[32] , 
        \R_DATA_TEMPR82[31] , \R_DATA_TEMPR82[30] , 
        \R_DATA_TEMPR82[29] , \R_DATA_TEMPR82[28] , 
        \R_DATA_TEMPR82[27] , \R_DATA_TEMPR82[26] , 
        \R_DATA_TEMPR82[25] , \R_DATA_TEMPR82[24] , 
        \R_DATA_TEMPR82[23] , \R_DATA_TEMPR82[22] , 
        \R_DATA_TEMPR82[21] , \R_DATA_TEMPR82[20] }), .B_DOUT({
        \R_DATA_TEMPR82[19] , \R_DATA_TEMPR82[18] , 
        \R_DATA_TEMPR82[17] , \R_DATA_TEMPR82[16] , 
        \R_DATA_TEMPR82[15] , \R_DATA_TEMPR82[14] , 
        \R_DATA_TEMPR82[13] , \R_DATA_TEMPR82[12] , 
        \R_DATA_TEMPR82[11] , \R_DATA_TEMPR82[10] , 
        \R_DATA_TEMPR82[9] , \R_DATA_TEMPR82[8] , \R_DATA_TEMPR82[7] , 
        \R_DATA_TEMPR82[6] , \R_DATA_TEMPR82[5] , \R_DATA_TEMPR82[4] , 
        \R_DATA_TEMPR82[3] , \R_DATA_TEMPR82[2] , \R_DATA_TEMPR82[1] , 
        \R_DATA_TEMPR82[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[82][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[20] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[20] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%53%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R53C0 (.A_DOUT({
        \R_DATA_TEMPR53[39] , \R_DATA_TEMPR53[38] , 
        \R_DATA_TEMPR53[37] , \R_DATA_TEMPR53[36] , 
        \R_DATA_TEMPR53[35] , \R_DATA_TEMPR53[34] , 
        \R_DATA_TEMPR53[33] , \R_DATA_TEMPR53[32] , 
        \R_DATA_TEMPR53[31] , \R_DATA_TEMPR53[30] , 
        \R_DATA_TEMPR53[29] , \R_DATA_TEMPR53[28] , 
        \R_DATA_TEMPR53[27] , \R_DATA_TEMPR53[26] , 
        \R_DATA_TEMPR53[25] , \R_DATA_TEMPR53[24] , 
        \R_DATA_TEMPR53[23] , \R_DATA_TEMPR53[22] , 
        \R_DATA_TEMPR53[21] , \R_DATA_TEMPR53[20] }), .B_DOUT({
        \R_DATA_TEMPR53[19] , \R_DATA_TEMPR53[18] , 
        \R_DATA_TEMPR53[17] , \R_DATA_TEMPR53[16] , 
        \R_DATA_TEMPR53[15] , \R_DATA_TEMPR53[14] , 
        \R_DATA_TEMPR53[13] , \R_DATA_TEMPR53[12] , 
        \R_DATA_TEMPR53[11] , \R_DATA_TEMPR53[10] , 
        \R_DATA_TEMPR53[9] , \R_DATA_TEMPR53[8] , \R_DATA_TEMPR53[7] , 
        \R_DATA_TEMPR53[6] , \R_DATA_TEMPR53[5] , \R_DATA_TEMPR53[4] , 
        \R_DATA_TEMPR53[3] , \R_DATA_TEMPR53[2] , \R_DATA_TEMPR53[1] , 
        \R_DATA_TEMPR53[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[53][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[13] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[13] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1018 (.A(OR4_955_Y), .B(OR4_179_Y), .C(OR4_974_Y), .D(
        OR4_1234_Y), .Y(OR4_1018_Y));
    OR4 OR4_65 (.A(\R_DATA_TEMPR0[17] ), .B(\R_DATA_TEMPR1[17] ), .C(
        \R_DATA_TEMPR2[17] ), .D(\R_DATA_TEMPR3[17] ), .Y(OR4_65_Y));
    OR4 OR4_1524 (.A(OR4_1333_Y), .B(OR4_1097_Y), .C(OR4_1080_Y), .D(
        OR4_761_Y), .Y(OR4_1524_Y));
    OR4 OR4_991 (.A(OR4_322_Y), .B(OR4_663_Y), .C(OR4_1200_Y), .D(
        OR4_603_Y), .Y(OR4_991_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%43%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R43C0 (.A_DOUT({
        \R_DATA_TEMPR43[39] , \R_DATA_TEMPR43[38] , 
        \R_DATA_TEMPR43[37] , \R_DATA_TEMPR43[36] , 
        \R_DATA_TEMPR43[35] , \R_DATA_TEMPR43[34] , 
        \R_DATA_TEMPR43[33] , \R_DATA_TEMPR43[32] , 
        \R_DATA_TEMPR43[31] , \R_DATA_TEMPR43[30] , 
        \R_DATA_TEMPR43[29] , \R_DATA_TEMPR43[28] , 
        \R_DATA_TEMPR43[27] , \R_DATA_TEMPR43[26] , 
        \R_DATA_TEMPR43[25] , \R_DATA_TEMPR43[24] , 
        \R_DATA_TEMPR43[23] , \R_DATA_TEMPR43[22] , 
        \R_DATA_TEMPR43[21] , \R_DATA_TEMPR43[20] }), .B_DOUT({
        \R_DATA_TEMPR43[19] , \R_DATA_TEMPR43[18] , 
        \R_DATA_TEMPR43[17] , \R_DATA_TEMPR43[16] , 
        \R_DATA_TEMPR43[15] , \R_DATA_TEMPR43[14] , 
        \R_DATA_TEMPR43[13] , \R_DATA_TEMPR43[12] , 
        \R_DATA_TEMPR43[11] , \R_DATA_TEMPR43[10] , 
        \R_DATA_TEMPR43[9] , \R_DATA_TEMPR43[8] , \R_DATA_TEMPR43[7] , 
        \R_DATA_TEMPR43[6] , \R_DATA_TEMPR43[5] , \R_DATA_TEMPR43[4] , 
        \R_DATA_TEMPR43[3] , \R_DATA_TEMPR43[2] , \R_DATA_TEMPR43[1] , 
        \R_DATA_TEMPR43[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[43][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[10] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[10] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_360 (.A(OR4_486_Y), .B(OR4_1393_Y), .C(OR4_386_Y), .D(
        OR4_1148_Y), .Y(OR4_360_Y));
    OR4 OR4_1325 (.A(\R_DATA_TEMPR68[39] ), .B(\R_DATA_TEMPR69[39] ), 
        .C(\R_DATA_TEMPR70[39] ), .D(\R_DATA_TEMPR71[39] ), .Y(
        OR4_1325_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%102%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R102C0 (.A_DOUT({
        \R_DATA_TEMPR102[39] , \R_DATA_TEMPR102[38] , 
        \R_DATA_TEMPR102[37] , \R_DATA_TEMPR102[36] , 
        \R_DATA_TEMPR102[35] , \R_DATA_TEMPR102[34] , 
        \R_DATA_TEMPR102[33] , \R_DATA_TEMPR102[32] , 
        \R_DATA_TEMPR102[31] , \R_DATA_TEMPR102[30] , 
        \R_DATA_TEMPR102[29] , \R_DATA_TEMPR102[28] , 
        \R_DATA_TEMPR102[27] , \R_DATA_TEMPR102[26] , 
        \R_DATA_TEMPR102[25] , \R_DATA_TEMPR102[24] , 
        \R_DATA_TEMPR102[23] , \R_DATA_TEMPR102[22] , 
        \R_DATA_TEMPR102[21] , \R_DATA_TEMPR102[20] }), .B_DOUT({
        \R_DATA_TEMPR102[19] , \R_DATA_TEMPR102[18] , 
        \R_DATA_TEMPR102[17] , \R_DATA_TEMPR102[16] , 
        \R_DATA_TEMPR102[15] , \R_DATA_TEMPR102[14] , 
        \R_DATA_TEMPR102[13] , \R_DATA_TEMPR102[12] , 
        \R_DATA_TEMPR102[11] , \R_DATA_TEMPR102[10] , 
        \R_DATA_TEMPR102[9] , \R_DATA_TEMPR102[8] , 
        \R_DATA_TEMPR102[7] , \R_DATA_TEMPR102[6] , 
        \R_DATA_TEMPR102[5] , \R_DATA_TEMPR102[4] , 
        \R_DATA_TEMPR102[3] , \R_DATA_TEMPR102[2] , 
        \R_DATA_TEMPR102[1] , \R_DATA_TEMPR102[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[102][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[25] , R_ADDR[10], \BLKY0[0] }), 
        .A_CLK(CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], 
        W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], 
        W_DATA[31], W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], 
        W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], 
        W_DATA[21], W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], 
        WBYTE_EN[2]}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], 
        W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], 
        W_ADDR[0], GND, GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[25] , 
        W_ADDR[10], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA[19], 
        W_DATA[18], W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], 
        W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], W_DATA[9], 
        W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], 
        W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_355 (.A(\R_DATA_TEMPR112[22] ), .B(\R_DATA_TEMPR113[22] ), 
        .C(\R_DATA_TEMPR114[22] ), .D(\R_DATA_TEMPR115[22] ), .Y(
        OR4_355_Y));
    OR4 OR4_1194 (.A(\R_DATA_TEMPR124[6] ), .B(\R_DATA_TEMPR125[6] ), 
        .C(\R_DATA_TEMPR126[6] ), .D(\R_DATA_TEMPR127[6] ), .Y(
        OR4_1194_Y));
    OR4 OR4_328 (.A(\R_DATA_TEMPR12[20] ), .B(\R_DATA_TEMPR13[20] ), 
        .C(\R_DATA_TEMPR14[20] ), .D(\R_DATA_TEMPR15[20] ), .Y(
        OR4_328_Y));
    OR4 OR4_344 (.A(\R_DATA_TEMPR108[30] ), .B(\R_DATA_TEMPR109[30] ), 
        .C(\R_DATA_TEMPR110[30] ), .D(\R_DATA_TEMPR111[30] ), .Y(
        OR4_344_Y));
    OR4 OR4_1512 (.A(OR4_814_Y), .B(OR4_359_Y), .C(OR4_339_Y), .D(
        OR4_1639_Y), .Y(OR4_1512_Y));
    OR4 OR4_863 (.A(\R_DATA_TEMPR80[6] ), .B(\R_DATA_TEMPR81[6] ), .C(
        \R_DATA_TEMPR82[6] ), .D(\R_DATA_TEMPR83[6] ), .Y(OR4_863_Y));
    OR4 OR4_185 (.A(\R_DATA_TEMPR8[16] ), .B(\R_DATA_TEMPR9[16] ), .C(
        \R_DATA_TEMPR10[16] ), .D(\R_DATA_TEMPR11[16] ), .Y(OR4_185_Y));
    OR4 OR4_1590 (.A(OR4_178_Y), .B(OR4_498_Y), .C(OR4_731_Y), .D(
        OR4_547_Y), .Y(OR4_1590_Y));
    OR4 OR4_141 (.A(\R_DATA_TEMPR108[8] ), .B(\R_DATA_TEMPR109[8] ), 
        .C(\R_DATA_TEMPR110[8] ), .D(\R_DATA_TEMPR111[8] ), .Y(
        OR4_141_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[16]  (.A(CFG3_16_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[16] ));
    OR4 OR4_717 (.A(OR4_1600_Y), .B(OR2_31_Y), .C(\R_DATA_TEMPR86[38] )
        , .D(\R_DATA_TEMPR87[38] ), .Y(OR4_717_Y));
    OR4 OR4_36 (.A(\R_DATA_TEMPR16[5] ), .B(\R_DATA_TEMPR17[5] ), .C(
        \R_DATA_TEMPR18[5] ), .D(\R_DATA_TEMPR19[5] ), .Y(OR4_36_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%5%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C0 (.A_DOUT({
        \R_DATA_TEMPR5[39] , \R_DATA_TEMPR5[38] , \R_DATA_TEMPR5[37] , 
        \R_DATA_TEMPR5[36] , \R_DATA_TEMPR5[35] , \R_DATA_TEMPR5[34] , 
        \R_DATA_TEMPR5[33] , \R_DATA_TEMPR5[32] , \R_DATA_TEMPR5[31] , 
        \R_DATA_TEMPR5[30] , \R_DATA_TEMPR5[29] , \R_DATA_TEMPR5[28] , 
        \R_DATA_TEMPR5[27] , \R_DATA_TEMPR5[26] , \R_DATA_TEMPR5[25] , 
        \R_DATA_TEMPR5[24] , \R_DATA_TEMPR5[23] , \R_DATA_TEMPR5[22] , 
        \R_DATA_TEMPR5[21] , \R_DATA_TEMPR5[20] }), .B_DOUT({
        \R_DATA_TEMPR5[19] , \R_DATA_TEMPR5[18] , \R_DATA_TEMPR5[17] , 
        \R_DATA_TEMPR5[16] , \R_DATA_TEMPR5[15] , \R_DATA_TEMPR5[14] , 
        \R_DATA_TEMPR5[13] , \R_DATA_TEMPR5[12] , \R_DATA_TEMPR5[11] , 
        \R_DATA_TEMPR5[10] , \R_DATA_TEMPR5[9] , \R_DATA_TEMPR5[8] , 
        \R_DATA_TEMPR5[7] , \R_DATA_TEMPR5[6] , \R_DATA_TEMPR5[5] , 
        \R_DATA_TEMPR5[4] , \R_DATA_TEMPR5[3] , \R_DATA_TEMPR5[2] , 
        \R_DATA_TEMPR5[1] , \R_DATA_TEMPR5[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[5][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1475 (.A(\R_DATA_TEMPR72[34] ), .B(\R_DATA_TEMPR73[34] ), 
        .C(\R_DATA_TEMPR74[34] ), .D(\R_DATA_TEMPR75[34] ), .Y(
        OR4_1475_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%61%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R61C0 (.A_DOUT({
        \R_DATA_TEMPR61[39] , \R_DATA_TEMPR61[38] , 
        \R_DATA_TEMPR61[37] , \R_DATA_TEMPR61[36] , 
        \R_DATA_TEMPR61[35] , \R_DATA_TEMPR61[34] , 
        \R_DATA_TEMPR61[33] , \R_DATA_TEMPR61[32] , 
        \R_DATA_TEMPR61[31] , \R_DATA_TEMPR61[30] , 
        \R_DATA_TEMPR61[29] , \R_DATA_TEMPR61[28] , 
        \R_DATA_TEMPR61[27] , \R_DATA_TEMPR61[26] , 
        \R_DATA_TEMPR61[25] , \R_DATA_TEMPR61[24] , 
        \R_DATA_TEMPR61[23] , \R_DATA_TEMPR61[22] , 
        \R_DATA_TEMPR61[21] , \R_DATA_TEMPR61[20] }), .B_DOUT({
        \R_DATA_TEMPR61[19] , \R_DATA_TEMPR61[18] , 
        \R_DATA_TEMPR61[17] , \R_DATA_TEMPR61[16] , 
        \R_DATA_TEMPR61[15] , \R_DATA_TEMPR61[14] , 
        \R_DATA_TEMPR61[13] , \R_DATA_TEMPR61[12] , 
        \R_DATA_TEMPR61[11] , \R_DATA_TEMPR61[10] , 
        \R_DATA_TEMPR61[9] , \R_DATA_TEMPR61[8] , \R_DATA_TEMPR61[7] , 
        \R_DATA_TEMPR61[6] , \R_DATA_TEMPR61[5] , \R_DATA_TEMPR61[4] , 
        \R_DATA_TEMPR61[3] , \R_DATA_TEMPR61[2] , \R_DATA_TEMPR61[1] , 
        \R_DATA_TEMPR61[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[61][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[15] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[15] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_487 (.A(\R_DATA_TEMPR0[0] ), .B(\R_DATA_TEMPR1[0] ), .C(
        \R_DATA_TEMPR2[0] ), .D(\R_DATA_TEMPR3[0] ), .Y(OR4_487_Y));
    OR4 OR4_714 (.A(\R_DATA_TEMPR24[21] ), .B(\R_DATA_TEMPR25[21] ), 
        .C(\R_DATA_TEMPR26[21] ), .D(\R_DATA_TEMPR27[21] ), .Y(
        OR4_714_Y));
    OR4 OR4_501 (.A(\R_DATA_TEMPR100[35] ), .B(\R_DATA_TEMPR101[35] ), 
        .C(\R_DATA_TEMPR102[35] ), .D(\R_DATA_TEMPR103[35] ), .Y(
        OR4_501_Y));
    CFG3 #( .INIT(8'h80) )  CFG3_23 (.A(W_ADDR[13]), .B(W_ADDR[12]), 
        .C(W_ADDR[11]), .Y(CFG3_23_Y));
    OR4 OR4_1555 (.A(\R_DATA_TEMPR116[14] ), .B(\R_DATA_TEMPR117[14] ), 
        .C(\R_DATA_TEMPR118[14] ), .D(\R_DATA_TEMPR119[14] ), .Y(
        OR4_1555_Y));
    OR4 OR4_21 (.A(\R_DATA_TEMPR120[37] ), .B(\R_DATA_TEMPR121[37] ), 
        .C(\R_DATA_TEMPR122[37] ), .D(\R_DATA_TEMPR123[37] ), .Y(
        OR4_21_Y));
    OR4 OR4_1298 (.A(\R_DATA_TEMPR16[15] ), .B(\R_DATA_TEMPR17[15] ), 
        .C(\R_DATA_TEMPR18[15] ), .D(\R_DATA_TEMPR19[15] ), .Y(
        OR4_1298_Y));
    OR4 OR4_1165 (.A(\R_DATA_TEMPR68[37] ), .B(\R_DATA_TEMPR69[37] ), 
        .C(\R_DATA_TEMPR70[37] ), .D(\R_DATA_TEMPR71[37] ), .Y(
        OR4_1165_Y));
    OR4 OR4_1107 (.A(\R_DATA_TEMPR24[34] ), .B(\R_DATA_TEMPR25[34] ), 
        .C(\R_DATA_TEMPR26[34] ), .D(\R_DATA_TEMPR27[34] ), .Y(
        OR4_1107_Y));
    OR4 OR4_937 (.A(OR4_794_Y), .B(OR4_543_Y), .C(OR4_258_Y), .D(
        OR4_1028_Y), .Y(OR4_937_Y));
    OR4 OR4_1032 (.A(OR4_1326_Y), .B(OR4_1627_Y), .C(OR4_1061_Y), .D(
        OR4_302_Y), .Y(OR4_1032_Y));
    OR4 OR4_129 (.A(\R_DATA_TEMPR24[24] ), .B(\R_DATA_TEMPR25[24] ), 
        .C(\R_DATA_TEMPR26[24] ), .D(\R_DATA_TEMPR27[24] ), .Y(
        OR4_129_Y));
    OR4 OR4_571 (.A(\R_DATA_TEMPR88[35] ), .B(\R_DATA_TEMPR89[35] ), 
        .C(\R_DATA_TEMPR90[35] ), .D(\R_DATA_TEMPR91[35] ), .Y(
        OR4_571_Y));
    OR4 OR4_1061 (.A(\R_DATA_TEMPR104[7] ), .B(\R_DATA_TEMPR105[7] ), 
        .C(\R_DATA_TEMPR106[7] ), .D(\R_DATA_TEMPR107[7] ), .Y(
        OR4_1061_Y));
    OR4 OR4_811 (.A(\R_DATA_TEMPR32[23] ), .B(\R_DATA_TEMPR33[23] ), 
        .C(\R_DATA_TEMPR34[23] ), .D(\R_DATA_TEMPR35[23] ), .Y(
        OR4_811_Y));
    OR4 OR4_1256 (.A(\R_DATA_TEMPR44[17] ), .B(\R_DATA_TEMPR45[17] ), 
        .C(\R_DATA_TEMPR46[17] ), .D(\R_DATA_TEMPR47[17] ), .Y(
        OR4_1256_Y));
    OR4 OR4_752 (.A(\R_DATA_TEMPR72[23] ), .B(\R_DATA_TEMPR73[23] ), 
        .C(\R_DATA_TEMPR74[23] ), .D(\R_DATA_TEMPR75[23] ), .Y(
        OR4_752_Y));
    OR4 OR4_441 (.A(OR4_130_Y), .B(OR4_489_Y), .C(OR4_1009_Y), .D(
        OR4_421_Y), .Y(OR4_441_Y));
    OR4 OR4_795 (.A(\R_DATA_TEMPR16[10] ), .B(\R_DATA_TEMPR17[10] ), 
        .C(\R_DATA_TEMPR18[10] ), .D(\R_DATA_TEMPR19[10] ), .Y(
        OR4_795_Y));
    OR4 OR4_697 (.A(\R_DATA_TEMPR32[15] ), .B(\R_DATA_TEMPR33[15] ), 
        .C(\R_DATA_TEMPR34[15] ), .D(\R_DATA_TEMPR35[15] ), .Y(
        OR4_697_Y));
    OR4 OR4_448 (.A(OR4_1164_Y), .B(OR4_1446_Y), .C(OR4_1629_Y), .D(
        OR4_842_Y), .Y(OR4_448_Y));
    OR4 OR4_796 (.A(\R_DATA_TEMPR92[37] ), .B(\R_DATA_TEMPR93[37] ), 
        .C(\R_DATA_TEMPR94[37] ), .D(\R_DATA_TEMPR95[37] ), .Y(
        OR4_796_Y));
    OR4 OR4_285 (.A(\R_DATA_TEMPR0[32] ), .B(\R_DATA_TEMPR1[32] ), .C(
        \R_DATA_TEMPR2[32] ), .D(\R_DATA_TEMPR3[32] ), .Y(OR4_285_Y));
    OR4 OR4_1358 (.A(OR4_404_Y), .B(OR4_657_Y), .C(OR4_846_Y), .D(
        OR4_1599_Y), .Y(OR4_1358_Y));
    OR4 OR4_956 (.A(\R_DATA_TEMPR120[6] ), .B(\R_DATA_TEMPR121[6] ), 
        .C(\R_DATA_TEMPR122[6] ), .D(\R_DATA_TEMPR123[6] ), .Y(
        OR4_956_Y));
    OR4 OR4_882 (.A(\R_DATA_TEMPR80[24] ), .B(\R_DATA_TEMPR81[24] ), 
        .C(\R_DATA_TEMPR82[24] ), .D(\R_DATA_TEMPR83[24] ), .Y(
        OR4_882_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%118%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R118C0 (.A_DOUT({
        \R_DATA_TEMPR118[39] , \R_DATA_TEMPR118[38] , 
        \R_DATA_TEMPR118[37] , \R_DATA_TEMPR118[36] , 
        \R_DATA_TEMPR118[35] , \R_DATA_TEMPR118[34] , 
        \R_DATA_TEMPR118[33] , \R_DATA_TEMPR118[32] , 
        \R_DATA_TEMPR118[31] , \R_DATA_TEMPR118[30] , 
        \R_DATA_TEMPR118[29] , \R_DATA_TEMPR118[28] , 
        \R_DATA_TEMPR118[27] , \R_DATA_TEMPR118[26] , 
        \R_DATA_TEMPR118[25] , \R_DATA_TEMPR118[24] , 
        \R_DATA_TEMPR118[23] , \R_DATA_TEMPR118[22] , 
        \R_DATA_TEMPR118[21] , \R_DATA_TEMPR118[20] }), .B_DOUT({
        \R_DATA_TEMPR118[19] , \R_DATA_TEMPR118[18] , 
        \R_DATA_TEMPR118[17] , \R_DATA_TEMPR118[16] , 
        \R_DATA_TEMPR118[15] , \R_DATA_TEMPR118[14] , 
        \R_DATA_TEMPR118[13] , \R_DATA_TEMPR118[12] , 
        \R_DATA_TEMPR118[11] , \R_DATA_TEMPR118[10] , 
        \R_DATA_TEMPR118[9] , \R_DATA_TEMPR118[8] , 
        \R_DATA_TEMPR118[7] , \R_DATA_TEMPR118[6] , 
        \R_DATA_TEMPR118[5] , \R_DATA_TEMPR118[4] , 
        \R_DATA_TEMPR118[3] , \R_DATA_TEMPR118[2] , 
        \R_DATA_TEMPR118[1] , \R_DATA_TEMPR118[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[118][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[29] , R_ADDR[10], \BLKY0[0] }), 
        .A_CLK(CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], 
        W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], 
        W_DATA[31], W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], 
        W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], 
        W_DATA[21], W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], 
        WBYTE_EN[2]}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], 
        W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], 
        W_ADDR[0], GND, GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[29] , 
        W_ADDR[10], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA[19], 
        W_DATA[18], W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], 
        W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], W_DATA[9], 
        W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], 
        W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_202 (.A(OR4_924_Y), .B(OR4_755_Y), .C(OR4_139_Y), .D(
        OR4_669_Y), .Y(OR4_202_Y));
    OR4 OR4_655 (.A(\R_DATA_TEMPR24[9] ), .B(\R_DATA_TEMPR25[9] ), .C(
        \R_DATA_TEMPR26[9] ), .D(\R_DATA_TEMPR27[9] ), .Y(OR4_655_Y));
    OR4 OR4_921 (.A(OR4_174_Y), .B(OR2_17_Y), .C(\R_DATA_TEMPR86[2] ), 
        .D(\R_DATA_TEMPR87[2] ), .Y(OR4_921_Y));
    OR4 OR4_1063 (.A(OR4_1397_Y), .B(OR4_209_Y), .C(OR4_1159_Y), .D(
        OR4_1489_Y), .Y(OR4_1063_Y));
    CFG3 #( .INIT(8'h1) )  CFG3_13 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_13_Y));
    OR4 OR4_272 (.A(\R_DATA_TEMPR16[39] ), .B(\R_DATA_TEMPR17[39] ), 
        .C(\R_DATA_TEMPR18[39] ), .D(\R_DATA_TEMPR19[39] ), .Y(
        OR4_272_Y));
    OR4 OR4_1462 (.A(\R_DATA_TEMPR72[25] ), .B(\R_DATA_TEMPR73[25] ), 
        .C(\R_DATA_TEMPR74[25] ), .D(\R_DATA_TEMPR75[25] ), .Y(
        OR4_1462_Y));
    OR4 OR4_1187 (.A(OR4_49_Y), .B(OR4_1178_Y), .C(OR4_1238_Y), .D(
        OR4_511_Y), .Y(OR4_1187_Y));
    OR4 OR4_1017 (.A(\R_DATA_TEMPR60[6] ), .B(\R_DATA_TEMPR61[6] ), .C(
        \R_DATA_TEMPR62[6] ), .D(\R_DATA_TEMPR63[6] ), .Y(OR4_1017_Y));
    OR4 OR4_1376 (.A(\R_DATA_TEMPR124[33] ), .B(\R_DATA_TEMPR125[33] ), 
        .C(\R_DATA_TEMPR126[33] ), .D(\R_DATA_TEMPR127[33] ), .Y(
        OR4_1376_Y));
    OR4 OR4_565 (.A(\R_DATA_TEMPR60[22] ), .B(\R_DATA_TEMPR61[22] ), 
        .C(\R_DATA_TEMPR62[22] ), .D(\R_DATA_TEMPR63[22] ), .Y(
        OR4_565_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%109%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R109C0 (.A_DOUT({
        \R_DATA_TEMPR109[39] , \R_DATA_TEMPR109[38] , 
        \R_DATA_TEMPR109[37] , \R_DATA_TEMPR109[36] , 
        \R_DATA_TEMPR109[35] , \R_DATA_TEMPR109[34] , 
        \R_DATA_TEMPR109[33] , \R_DATA_TEMPR109[32] , 
        \R_DATA_TEMPR109[31] , \R_DATA_TEMPR109[30] , 
        \R_DATA_TEMPR109[29] , \R_DATA_TEMPR109[28] , 
        \R_DATA_TEMPR109[27] , \R_DATA_TEMPR109[26] , 
        \R_DATA_TEMPR109[25] , \R_DATA_TEMPR109[24] , 
        \R_DATA_TEMPR109[23] , \R_DATA_TEMPR109[22] , 
        \R_DATA_TEMPR109[21] , \R_DATA_TEMPR109[20] }), .B_DOUT({
        \R_DATA_TEMPR109[19] , \R_DATA_TEMPR109[18] , 
        \R_DATA_TEMPR109[17] , \R_DATA_TEMPR109[16] , 
        \R_DATA_TEMPR109[15] , \R_DATA_TEMPR109[14] , 
        \R_DATA_TEMPR109[13] , \R_DATA_TEMPR109[12] , 
        \R_DATA_TEMPR109[11] , \R_DATA_TEMPR109[10] , 
        \R_DATA_TEMPR109[9] , \R_DATA_TEMPR109[8] , 
        \R_DATA_TEMPR109[7] , \R_DATA_TEMPR109[6] , 
        \R_DATA_TEMPR109[5] , \R_DATA_TEMPR109[4] , 
        \R_DATA_TEMPR109[3] , \R_DATA_TEMPR109[2] , 
        \R_DATA_TEMPR109[1] , \R_DATA_TEMPR109[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[109][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[27] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[27] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_44 (.A(\R_DATA_TEMPR40[32] ), .B(\R_DATA_TEMPR41[32] ), .C(
        \R_DATA_TEMPR42[32] ), .D(\R_DATA_TEMPR43[32] ), .Y(OR4_44_Y));
    OR4 OR4_549 (.A(\R_DATA_TEMPR80[39] ), .B(\R_DATA_TEMPR81[39] ), 
        .C(\R_DATA_TEMPR82[39] ), .D(\R_DATA_TEMPR83[39] ), .Y(
        OR4_549_Y));
    OR4 OR4_300 (.A(\R_DATA_TEMPR24[27] ), .B(\R_DATA_TEMPR25[27] ), 
        .C(\R_DATA_TEMPR26[27] ), .D(\R_DATA_TEMPR27[27] ), .Y(
        OR4_300_Y));
    OR4 OR4_435 (.A(\R_DATA_TEMPR16[18] ), .B(\R_DATA_TEMPR17[18] ), 
        .C(\R_DATA_TEMPR18[18] ), .D(\R_DATA_TEMPR19[18] ), .Y(
        OR4_435_Y));
    OR4 OR4_540 (.A(\R_DATA_TEMPR40[23] ), .B(\R_DATA_TEMPR41[23] ), 
        .C(\R_DATA_TEMPR42[23] ), .D(\R_DATA_TEMPR43[23] ), .Y(
        OR4_540_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%91%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R91C0 (.A_DOUT({
        \R_DATA_TEMPR91[39] , \R_DATA_TEMPR91[38] , 
        \R_DATA_TEMPR91[37] , \R_DATA_TEMPR91[36] , 
        \R_DATA_TEMPR91[35] , \R_DATA_TEMPR91[34] , 
        \R_DATA_TEMPR91[33] , \R_DATA_TEMPR91[32] , 
        \R_DATA_TEMPR91[31] , \R_DATA_TEMPR91[30] , 
        \R_DATA_TEMPR91[29] , \R_DATA_TEMPR91[28] , 
        \R_DATA_TEMPR91[27] , \R_DATA_TEMPR91[26] , 
        \R_DATA_TEMPR91[25] , \R_DATA_TEMPR91[24] , 
        \R_DATA_TEMPR91[23] , \R_DATA_TEMPR91[22] , 
        \R_DATA_TEMPR91[21] , \R_DATA_TEMPR91[20] }), .B_DOUT({
        \R_DATA_TEMPR91[19] , \R_DATA_TEMPR91[18] , 
        \R_DATA_TEMPR91[17] , \R_DATA_TEMPR91[16] , 
        \R_DATA_TEMPR91[15] , \R_DATA_TEMPR91[14] , 
        \R_DATA_TEMPR91[13] , \R_DATA_TEMPR91[12] , 
        \R_DATA_TEMPR91[11] , \R_DATA_TEMPR91[10] , 
        \R_DATA_TEMPR91[9] , \R_DATA_TEMPR91[8] , \R_DATA_TEMPR91[7] , 
        \R_DATA_TEMPR91[6] , \R_DATA_TEMPR91[5] , \R_DATA_TEMPR91[4] , 
        \R_DATA_TEMPR91[3] , \R_DATA_TEMPR91[2] , \R_DATA_TEMPR91[1] , 
        \R_DATA_TEMPR91[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[91][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[22] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[22] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_483 (.A(\R_DATA_TEMPR80[23] ), .B(\R_DATA_TEMPR81[23] ), 
        .C(\R_DATA_TEMPR82[23] ), .D(\R_DATA_TEMPR83[23] ), .Y(
        OR4_483_Y));
    OR4 OR4_1243 (.A(OR4_1604_Y), .B(OR4_224_Y), .C(OR4_1370_Y), .D(
        OR4_1094_Y), .Y(OR4_1243_Y));
    OR4 OR4_1059 (.A(OR4_1084_Y), .B(OR4_26_Y), .C(OR4_815_Y), .D(
        OR4_1067_Y), .Y(OR4_1059_Y));
    OR4 OR4_681 (.A(\R_DATA_TEMPR36[25] ), .B(\R_DATA_TEMPR37[25] ), 
        .C(\R_DATA_TEMPR38[25] ), .D(\R_DATA_TEMPR39[25] ), .Y(
        OR4_681_Y));
    OR4 OR4_663 (.A(OR4_198_Y), .B(OR2_29_Y), .C(\R_DATA_TEMPR86[22] ), 
        .D(\R_DATA_TEMPR87[22] ), .Y(OR4_663_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[22]  (.A(CFG3_1_Y), .B(CFG3_9_Y)
        , .Y(\BLKY2[22] ));
    OR4 OR4_1195 (.A(OR4_1064_Y), .B(OR4_727_Y), .C(OR4_1085_Y), .D(
        OR4_197_Y), .Y(OR4_1195_Y));
    OR4 OR4_370 (.A(\R_DATA_TEMPR64[25] ), .B(\R_DATA_TEMPR65[25] ), 
        .C(\R_DATA_TEMPR66[25] ), .D(\R_DATA_TEMPR67[25] ), .Y(
        OR4_370_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%6%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C0 (.A_DOUT({
        \R_DATA_TEMPR6[39] , \R_DATA_TEMPR6[38] , \R_DATA_TEMPR6[37] , 
        \R_DATA_TEMPR6[36] , \R_DATA_TEMPR6[35] , \R_DATA_TEMPR6[34] , 
        \R_DATA_TEMPR6[33] , \R_DATA_TEMPR6[32] , \R_DATA_TEMPR6[31] , 
        \R_DATA_TEMPR6[30] , \R_DATA_TEMPR6[29] , \R_DATA_TEMPR6[28] , 
        \R_DATA_TEMPR6[27] , \R_DATA_TEMPR6[26] , \R_DATA_TEMPR6[25] , 
        \R_DATA_TEMPR6[24] , \R_DATA_TEMPR6[23] , \R_DATA_TEMPR6[22] , 
        \R_DATA_TEMPR6[21] , \R_DATA_TEMPR6[20] }), .B_DOUT({
        \R_DATA_TEMPR6[19] , \R_DATA_TEMPR6[18] , \R_DATA_TEMPR6[17] , 
        \R_DATA_TEMPR6[16] , \R_DATA_TEMPR6[15] , \R_DATA_TEMPR6[14] , 
        \R_DATA_TEMPR6[13] , \R_DATA_TEMPR6[12] , \R_DATA_TEMPR6[11] , 
        \R_DATA_TEMPR6[10] , \R_DATA_TEMPR6[9] , \R_DATA_TEMPR6[8] , 
        \R_DATA_TEMPR6[7] , \R_DATA_TEMPR6[6] , \R_DATA_TEMPR6[5] , 
        \R_DATA_TEMPR6[4] , \R_DATA_TEMPR6[3] , \R_DATA_TEMPR6[2] , 
        \R_DATA_TEMPR6[1] , \R_DATA_TEMPR6[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[6][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_288 (.A(\R_DATA_TEMPR8[5] ), .B(\R_DATA_TEMPR9[5] ), .C(
        \R_DATA_TEMPR10[5] ), .D(\R_DATA_TEMPR11[5] ), .Y(OR4_288_Y));
    OR4 OR4_917 (.A(OR4_1369_Y), .B(OR4_756_Y), .C(OR4_994_Y), .D(
        OR4_1583_Y), .Y(OR4_917_Y));
    CFG3 #( .INIT(8'h4) )  CFG3_0 (.A(R_ADDR[13]), .B(R_ADDR[12]), .C(
        R_ADDR[11]), .Y(CFG3_0_Y));
    OR4 OR4_1022 (.A(\R_DATA_TEMPR64[32] ), .B(\R_DATA_TEMPR65[32] ), 
        .C(\R_DATA_TEMPR66[32] ), .D(\R_DATA_TEMPR67[32] ), .Y(
        OR4_1022_Y));
    OR4 OR4_1091 (.A(\R_DATA_TEMPR64[26] ), .B(\R_DATA_TEMPR65[26] ), 
        .C(\R_DATA_TEMPR66[26] ), .D(\R_DATA_TEMPR67[26] ), .Y(
        OR4_1091_Y));
    OR4 OR4_803 (.A(OR4_1348_Y), .B(OR4_1013_Y), .C(OR4_1467_Y), .D(
        OR4_1273_Y), .Y(OR4_803_Y));
    OR4 OR4_1200 (.A(\R_DATA_TEMPR88[22] ), .B(\R_DATA_TEMPR89[22] ), 
        .C(\R_DATA_TEMPR90[22] ), .D(\R_DATA_TEMPR91[22] ), .Y(
        OR4_1200_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[8]  (.A(CFG3_16_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[8] ));
    OR4 OR4_1533 (.A(\R_DATA_TEMPR120[7] ), .B(\R_DATA_TEMPR121[7] ), 
        .C(\R_DATA_TEMPR122[7] ), .D(\R_DATA_TEMPR123[7] ), .Y(
        OR4_1533_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[12]  (.A(CFG3_6_Y), .B(CFG3_4_Y)
        , .Y(\BLKX2[12] ));
    OR4 OR4_30 (.A(\R_DATA_TEMPR20[17] ), .B(\R_DATA_TEMPR21[17] ), .C(
        \R_DATA_TEMPR22[17] ), .D(\R_DATA_TEMPR23[17] ), .Y(OR4_30_Y));
    OR4 OR4_650 (.A(\R_DATA_TEMPR104[18] ), .B(\R_DATA_TEMPR105[18] ), 
        .C(\R_DATA_TEMPR106[18] ), .D(\R_DATA_TEMPR107[18] ), .Y(
        OR4_650_Y));
    OR4 OR4_873 (.A(\R_DATA_TEMPR12[39] ), .B(\R_DATA_TEMPR13[39] ), 
        .C(\R_DATA_TEMPR14[39] ), .D(\R_DATA_TEMPR15[39] ), .Y(
        OR4_873_Y));
    OR4 OR4_725 (.A(\R_DATA_TEMPR52[6] ), .B(\R_DATA_TEMPR53[6] ), .C(
        \R_DATA_TEMPR54[6] ), .D(\R_DATA_TEMPR55[6] ), .Y(OR4_725_Y));
    OR4 OR4_627 (.A(\R_DATA_TEMPR116[33] ), .B(\R_DATA_TEMPR117[33] ), 
        .C(\R_DATA_TEMPR118[33] ), .D(\R_DATA_TEMPR119[33] ), .Y(
        OR4_627_Y));
    OR4 OR4_297 (.A(OR4_1226_Y), .B(OR4_1044_Y), .C(OR4_453_Y), .D(
        OR4_968_Y), .Y(OR4_297_Y));
    OR4 OR4_1618 (.A(\R_DATA_TEMPR76[38] ), .B(\R_DATA_TEMPR77[38] ), 
        .C(\R_DATA_TEMPR78[38] ), .D(\R_DATA_TEMPR79[38] ), .Y(
        OR4_1618_Y));
    OR4 OR4_726 (.A(\R_DATA_TEMPR0[19] ), .B(\R_DATA_TEMPR1[19] ), .C(
        \R_DATA_TEMPR2[19] ), .D(\R_DATA_TEMPR3[19] ), .Y(OR4_726_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%0%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C0 (.A_DOUT({
        \R_DATA_TEMPR0[39] , \R_DATA_TEMPR0[38] , \R_DATA_TEMPR0[37] , 
        \R_DATA_TEMPR0[36] , \R_DATA_TEMPR0[35] , \R_DATA_TEMPR0[34] , 
        \R_DATA_TEMPR0[33] , \R_DATA_TEMPR0[32] , \R_DATA_TEMPR0[31] , 
        \R_DATA_TEMPR0[30] , \R_DATA_TEMPR0[29] , \R_DATA_TEMPR0[28] , 
        \R_DATA_TEMPR0[27] , \R_DATA_TEMPR0[26] , \R_DATA_TEMPR0[25] , 
        \R_DATA_TEMPR0[24] , \R_DATA_TEMPR0[23] , \R_DATA_TEMPR0[22] , 
        \R_DATA_TEMPR0[21] , \R_DATA_TEMPR0[20] }), .B_DOUT({
        \R_DATA_TEMPR0[19] , \R_DATA_TEMPR0[18] , \R_DATA_TEMPR0[17] , 
        \R_DATA_TEMPR0[16] , \R_DATA_TEMPR0[15] , \R_DATA_TEMPR0[14] , 
        \R_DATA_TEMPR0[13] , \R_DATA_TEMPR0[12] , \R_DATA_TEMPR0[11] , 
        \R_DATA_TEMPR0[10] , \R_DATA_TEMPR0[9] , \R_DATA_TEMPR0[8] , 
        \R_DATA_TEMPR0[7] , \R_DATA_TEMPR0[6] , \R_DATA_TEMPR0[5] , 
        \R_DATA_TEMPR0[4] , \R_DATA_TEMPR0[3] , \R_DATA_TEMPR0[2] , 
        \R_DATA_TEMPR0[1] , \R_DATA_TEMPR0[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[0][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1507 (.A(\R_DATA_TEMPR112[10] ), .B(\R_DATA_TEMPR113[10] ), 
        .C(\R_DATA_TEMPR114[10] ), .D(\R_DATA_TEMPR115[10] ), .Y(
        OR4_1507_Y));
    OR4 OR4_37 (.A(\R_DATA_TEMPR0[26] ), .B(\R_DATA_TEMPR1[26] ), .C(
        \R_DATA_TEMPR2[26] ), .D(\R_DATA_TEMPR3[26] ), .Y(OR4_37_Y));
    OR4 OR4_969 (.A(\R_DATA_TEMPR92[24] ), .B(\R_DATA_TEMPR93[24] ), 
        .C(\R_DATA_TEMPR94[24] ), .D(\R_DATA_TEMPR95[24] ), .Y(
        OR4_969_Y));
    OR4 OR4_960 (.A(OR4_1251_Y), .B(OR4_194_Y), .C(OR4_975_Y), .D(
        OR4_1237_Y), .Y(OR4_960_Y));
    OR4 OR4_197 (.A(OR4_484_Y), .B(OR4_1050_Y), .C(OR4_214_Y), .D(
        OR4_471_Y), .Y(OR4_197_Y));
    OR4 OR4_1302 (.A(\R_DATA_TEMPR108[16] ), .B(\R_DATA_TEMPR109[16] ), 
        .C(\R_DATA_TEMPR110[16] ), .D(\R_DATA_TEMPR111[16] ), .Y(
        OR4_1302_Y));
    OR4 OR4_1149 (.A(\R_DATA_TEMPR124[15] ), .B(\R_DATA_TEMPR125[15] ), 
        .C(\R_DATA_TEMPR126[15] ), .D(\R_DATA_TEMPR127[15] ), .Y(
        OR4_1149_Y));
    OR4 OR4_1478 (.A(\R_DATA_TEMPR112[30] ), .B(\R_DATA_TEMPR113[30] ), 
        .C(\R_DATA_TEMPR114[30] ), .D(\R_DATA_TEMPR115[30] ), .Y(
        OR4_1478_Y));
    OR4 OR4_1093 (.A(\R_DATA_TEMPR44[29] ), .B(\R_DATA_TEMPR45[29] ), 
        .C(\R_DATA_TEMPR46[29] ), .D(\R_DATA_TEMPR47[29] ), .Y(
        OR4_1093_Y));
    OR4 OR4_357 (.A(\R_DATA_TEMPR40[35] ), .B(\R_DATA_TEMPR41[35] ), 
        .C(\R_DATA_TEMPR42[35] ), .D(\R_DATA_TEMPR43[35] ), .Y(
        OR4_357_Y));
    OR4 OR4_150 (.A(OR4_280_Y), .B(OR4_1420_Y), .C(OR4_1475_Y), .D(
        OR4_14_Y), .Y(OR4_150_Y));
    OR4 OR4_434 (.A(\R_DATA_TEMPR16[4] ), .B(\R_DATA_TEMPR17[4] ), .C(
        \R_DATA_TEMPR18[4] ), .D(\R_DATA_TEMPR19[4] ), .Y(OR4_434_Y));
    OR4 OR4_1202 (.A(\R_DATA_TEMPR108[24] ), .B(\R_DATA_TEMPR109[24] ), 
        .C(\R_DATA_TEMPR110[24] ), .D(\R_DATA_TEMPR111[24] ), .Y(
        OR4_1202_Y));
    OR4 OR4_1492 (.A(\R_DATA_TEMPR100[8] ), .B(\R_DATA_TEMPR101[8] ), 
        .C(\R_DATA_TEMPR102[8] ), .D(\R_DATA_TEMPR103[8] ), .Y(
        OR4_1492_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[26]  (.A(CFG3_14_Y), .B(
        CFG3_7_Y), .Y(\BLKX2[26] ));
    CFG3 #( .INIT(8'h20) )  CFG3_20 (.A(R_EN), .B(R_ADDR[15]), .C(
        R_ADDR[14]), .Y(CFG3_20_Y));
    OR4 OR4_163 (.A(OR4_429_Y), .B(OR4_996_Y), .C(OR4_145_Y), .D(
        OR4_420_Y), .Y(OR4_163_Y));
    OR4 OR4_1068 (.A(\R_DATA_TEMPR52[18] ), .B(\R_DATA_TEMPR53[18] ), 
        .C(\R_DATA_TEMPR54[18] ), .D(\R_DATA_TEMPR55[18] ), .Y(
        OR4_1068_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%13%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C0 (.A_DOUT({
        \R_DATA_TEMPR13[39] , \R_DATA_TEMPR13[38] , 
        \R_DATA_TEMPR13[37] , \R_DATA_TEMPR13[36] , 
        \R_DATA_TEMPR13[35] , \R_DATA_TEMPR13[34] , 
        \R_DATA_TEMPR13[33] , \R_DATA_TEMPR13[32] , 
        \R_DATA_TEMPR13[31] , \R_DATA_TEMPR13[30] , 
        \R_DATA_TEMPR13[29] , \R_DATA_TEMPR13[28] , 
        \R_DATA_TEMPR13[27] , \R_DATA_TEMPR13[26] , 
        \R_DATA_TEMPR13[25] , \R_DATA_TEMPR13[24] , 
        \R_DATA_TEMPR13[23] , \R_DATA_TEMPR13[22] , 
        \R_DATA_TEMPR13[21] , \R_DATA_TEMPR13[20] }), .B_DOUT({
        \R_DATA_TEMPR13[19] , \R_DATA_TEMPR13[18] , 
        \R_DATA_TEMPR13[17] , \R_DATA_TEMPR13[16] , 
        \R_DATA_TEMPR13[15] , \R_DATA_TEMPR13[14] , 
        \R_DATA_TEMPR13[13] , \R_DATA_TEMPR13[12] , 
        \R_DATA_TEMPR13[11] , \R_DATA_TEMPR13[10] , 
        \R_DATA_TEMPR13[9] , \R_DATA_TEMPR13[8] , \R_DATA_TEMPR13[7] , 
        \R_DATA_TEMPR13[6] , \R_DATA_TEMPR13[5] , \R_DATA_TEMPR13[4] , 
        \R_DATA_TEMPR13[3] , \R_DATA_TEMPR13[2] , \R_DATA_TEMPR13[1] , 
        \R_DATA_TEMPR13[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_758 (.A(OR4_812_Y), .B(OR4_708_Y), .C(OR4_684_Y), .D(
        OR4_374_Y), .Y(OR4_758_Y));
    OR4 OR4_343 (.A(OR4_961_Y), .B(OR4_1271_Y), .C(OR4_723_Y), .D(
        OR4_1577_Y), .Y(OR4_343_Y));
    OR4 OR4_740 (.A(\R_DATA_TEMPR64[8] ), .B(\R_DATA_TEMPR65[8] ), .C(
        \R_DATA_TEMPR66[8] ), .D(\R_DATA_TEMPR67[8] ), .Y(OR4_740_Y));
    OR4 OR4_336 (.A(\R_DATA_TEMPR44[22] ), .B(\R_DATA_TEMPR45[22] ), 
        .C(\R_DATA_TEMPR46[22] ), .D(\R_DATA_TEMPR47[22] ), .Y(
        OR4_336_Y));
    OR4 OR4_1404 (.A(\R_DATA_TEMPR32[30] ), .B(\R_DATA_TEMPR33[30] ), 
        .C(\R_DATA_TEMPR34[30] ), .D(\R_DATA_TEMPR35[30] ), .Y(
        OR4_1404_Y));
    OR4 OR4_1280 (.A(OR4_15_Y), .B(OR4_880_Y), .C(OR4_39_Y), .D(
        OR4_318_Y), .Y(OR4_1280_Y));
    OR4 OR4_415 (.A(\R_DATA_TEMPR12[11] ), .B(\R_DATA_TEMPR13[11] ), 
        .C(\R_DATA_TEMPR14[11] ), .D(\R_DATA_TEMPR15[11] ), .Y(
        OR4_415_Y));
    OR4 OR4_793 (.A(\R_DATA_TEMPR8[22] ), .B(\R_DATA_TEMPR9[22] ), .C(
        \R_DATA_TEMPR10[22] ), .D(\R_DATA_TEMPR11[22] ), .Y(OR4_793_Y));
    OR4 OR4_442 (.A(\R_DATA_TEMPR72[16] ), .B(\R_DATA_TEMPR73[16] ), 
        .C(\R_DATA_TEMPR74[16] ), .D(\R_DATA_TEMPR75[16] ), .Y(
        OR4_442_Y));
    OR4 OR4_1204 (.A(\R_DATA_TEMPR108[28] ), .B(\R_DATA_TEMPR109[28] ), 
        .C(\R_DATA_TEMPR110[28] ), .D(\R_DATA_TEMPR111[28] ), .Y(
        OR4_1204_Y));
    OR4 OR4_294 (.A(\R_DATA_TEMPR88[0] ), .B(\R_DATA_TEMPR89[0] ), .C(
        \R_DATA_TEMPR90[0] ), .D(\R_DATA_TEMPR91[0] ), .Y(OR4_294_Y));
    OR4 OR4_1562 (.A(\R_DATA_TEMPR88[13] ), .B(\R_DATA_TEMPR89[13] ), 
        .C(\R_DATA_TEMPR90[13] ), .D(\R_DATA_TEMPR91[13] ), .Y(
        OR4_1562_Y));
    OR4 OR4_1587 (.A(OR4_853_Y), .B(OR4_538_Y), .C(OR4_952_Y), .D(
        OR4_778_Y), .Y(OR4_1587_Y));
    OR4 OR4_449 (.A(\R_DATA_TEMPR120[36] ), .B(\R_DATA_TEMPR121[36] ), 
        .C(\R_DATA_TEMPR122[36] ), .D(\R_DATA_TEMPR123[36] ), .Y(
        OR4_449_Y));
    OR4 OR4_1174 (.A(\R_DATA_TEMPR12[9] ), .B(\R_DATA_TEMPR13[9] ), .C(
        \R_DATA_TEMPR14[9] ), .D(\R_DATA_TEMPR15[9] ), .Y(OR4_1174_Y));
    OR4 OR4_505 (.A(\R_DATA_TEMPR24[28] ), .B(\R_DATA_TEMPR25[28] ), 
        .C(\R_DATA_TEMPR26[28] ), .D(\R_DATA_TEMPR27[28] ), .Y(
        OR4_505_Y));
    OR4 OR4_1307 (.A(\R_DATA_TEMPR52[10] ), .B(\R_DATA_TEMPR53[10] ), 
        .C(\R_DATA_TEMPR54[10] ), .D(\R_DATA_TEMPR55[10] ), .Y(
        OR4_1307_Y));
    OR4 \OR4_R_DATA[24]  (.A(OR4_1428_Y), .B(OR4_851_Y), .C(OR4_8_Y), 
        .D(OR4_722_Y), .Y(R_DATA[24]));
    OR4 OR4_85 (.A(OR4_855_Y), .B(OR4_717_Y), .C(OR4_693_Y), .D(
        OR4_380_Y), .Y(OR4_85_Y));
    OR4 OR4_1382 (.A(\R_DATA_TEMPR76[0] ), .B(\R_DATA_TEMPR77[0] ), .C(
        \R_DATA_TEMPR78[0] ), .D(\R_DATA_TEMPR79[0] ), .Y(OR4_1382_Y));
    OR4 OR4_857 (.A(\R_DATA_TEMPR52[34] ), .B(\R_DATA_TEMPR53[34] ), 
        .C(\R_DATA_TEMPR54[34] ), .D(\R_DATA_TEMPR55[34] ), .Y(
        OR4_857_Y));
    OR4 OR4_146 (.A(\R_DATA_TEMPR80[8] ), .B(\R_DATA_TEMPR81[8] ), .C(
        \R_DATA_TEMPR82[8] ), .D(\R_DATA_TEMPR83[8] ), .Y(OR4_146_Y));
    OR4 OR4_158 (.A(OR4_803_Y), .B(OR4_115_Y), .C(OR4_188_Y), .D(
        OR4_1011_Y), .Y(OR4_158_Y));
    OR4 \OR4_R_DATA[12]  (.A(OR4_1171_Y), .B(OR4_1128_Y), .C(OR4_907_Y)
        , .D(OR4_170_Y), .Y(R_DATA[12]));
    OR4 OR4_954 (.A(\R_DATA_TEMPR124[39] ), .B(\R_DATA_TEMPR125[39] ), 
        .C(\R_DATA_TEMPR126[39] ), .D(\R_DATA_TEMPR127[39] ), .Y(
        OR4_954_Y));
    OR4 OR4_1523 (.A(OR4_819_Y), .B(OR4_71_Y), .C(OR4_44_Y), .D(
        OR4_1368_Y), .Y(OR4_1523_Y));
    OR4 OR4_1282 (.A(OR4_933_Y), .B(OR4_672_Y), .C(OR4_399_Y), .D(
        OR4_353_Y), .Y(OR4_1282_Y));
    OR4 OR4_1146 (.A(\R_DATA_TEMPR56[7] ), .B(\R_DATA_TEMPR57[7] ), .C(
        \R_DATA_TEMPR58[7] ), .D(\R_DATA_TEMPR59[7] ), .Y(OR4_1146_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_10 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_10_Y));
    OR4 OR4_1570 (.A(\R_DATA_TEMPR68[36] ), .B(\R_DATA_TEMPR69[36] ), 
        .C(\R_DATA_TEMPR70[36] ), .D(\R_DATA_TEMPR71[36] ), .Y(
        OR4_1570_Y));
    OR4 OR4_1441 (.A(OR4_370_Y), .B(OR4_104_Y), .C(OR4_1462_Y), .D(
        OR4_226_Y), .Y(OR4_1441_Y));
    OR4 OR4_581 (.A(\R_DATA_TEMPR0[16] ), .B(\R_DATA_TEMPR1[16] ), .C(
        \R_DATA_TEMPR2[16] ), .D(\R_DATA_TEMPR3[16] ), .Y(OR4_581_Y));
    OR4 OR4_575 (.A(\R_DATA_TEMPR88[11] ), .B(\R_DATA_TEMPR89[11] ), 
        .C(\R_DATA_TEMPR90[11] ), .D(\R_DATA_TEMPR91[11] ), .Y(
        OR4_575_Y));
    OR4 OR4_603 (.A(\R_DATA_TEMPR92[22] ), .B(\R_DATA_TEMPR93[22] ), 
        .C(\R_DATA_TEMPR94[22] ), .D(\R_DATA_TEMPR95[22] ), .Y(
        OR4_603_Y));
    OR4 OR4_69 (.A(\R_DATA_TEMPR0[12] ), .B(\R_DATA_TEMPR1[12] ), .C(
        \R_DATA_TEMPR2[12] ), .D(\R_DATA_TEMPR3[12] ), .Y(OR4_69_Y));
    OR4 OR4_1241 (.A(\R_DATA_TEMPR32[31] ), .B(\R_DATA_TEMPR33[31] ), 
        .C(\R_DATA_TEMPR34[31] ), .D(\R_DATA_TEMPR35[31] ), .Y(
        OR4_1241_Y));
    OR4 OR4_1615 (.A(\R_DATA_TEMPR116[37] ), .B(\R_DATA_TEMPR117[37] ), 
        .C(\R_DATA_TEMPR118[37] ), .D(\R_DATA_TEMPR119[37] ), .Y(
        OR4_1615_Y));
    OR4 OR4_1148 (.A(OR4_92_Y), .B(OR4_406_Y), .C(OR4_641_Y), .D(
        OR4_452_Y), .Y(OR4_1148_Y));
    OR4 OR4_1484 (.A(\R_DATA_TEMPR100[36] ), .B(\R_DATA_TEMPR101[36] ), 
        .C(\R_DATA_TEMPR102[36] ), .D(\R_DATA_TEMPR103[36] ), .Y(
        OR4_1484_Y));
    OR4 OR4_1157 (.A(\R_DATA_TEMPR36[29] ), .B(\R_DATA_TEMPR37[29] ), 
        .C(\R_DATA_TEMPR38[29] ), .D(\R_DATA_TEMPR39[29] ), .Y(
        OR4_1157_Y));
    OR4 OR4_227 (.A(\R_DATA_TEMPR48[19] ), .B(\R_DATA_TEMPR49[19] ), 
        .C(\R_DATA_TEMPR50[19] ), .D(\R_DATA_TEMPR51[19] ), .Y(
        OR4_227_Y));
    OR4 OR4_1278 (.A(\R_DATA_TEMPR16[6] ), .B(\R_DATA_TEMPR17[6] ), .C(
        \R_DATA_TEMPR18[6] ), .D(\R_DATA_TEMPR19[6] ), .Y(OR4_1278_Y));
    OR4 OR4_673 (.A(\R_DATA_TEMPR64[13] ), .B(\R_DATA_TEMPR65[13] ), 
        .C(\R_DATA_TEMPR66[13] ), .D(\R_DATA_TEMPR67[13] ), .Y(
        OR4_673_Y));
    OR4 OR4_1217 (.A(\R_DATA_TEMPR92[36] ), .B(\R_DATA_TEMPR93[36] ), 
        .C(\R_DATA_TEMPR94[36] ), .D(\R_DATA_TEMPR95[36] ), .Y(
        OR4_1217_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[21]  (.A(CFG3_11_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[21] ));
    OR4 OR4_395 (.A(OR4_926_Y), .B(OR4_770_Y), .C(OR4_896_Y), .D(
        OR4_607_Y), .Y(OR4_395_Y));
    OR4 OR4_414 (.A(\R_DATA_TEMPR44[31] ), .B(\R_DATA_TEMPR45[31] ), 
        .C(\R_DATA_TEMPR46[31] ), .D(\R_DATA_TEMPR47[31] ), .Y(
        OR4_414_Y));
    OR4 OR4_127 (.A(OR4_732_Y), .B(OR2_37_Y), .C(\R_DATA_TEMPR86[12] ), 
        .D(\R_DATA_TEMPR87[12] ), .Y(OR4_127_Y));
    OR4 OR4_1284 (.A(\R_DATA_TEMPR116[2] ), .B(\R_DATA_TEMPR117[2] ), 
        .C(\R_DATA_TEMPR118[2] ), .D(\R_DATA_TEMPR119[2] ), .Y(
        OR4_1284_Y));
    OR4 OR4_860 (.A(OR4_277_Y), .B(OR4_1593_Y), .C(OR4_384_Y), .D(
        OR4_211_Y), .Y(OR4_860_Y));
    OR4 OR4_348 (.A(OR4_983_Y), .B(OR4_1307_Y), .C(OR4_1538_Y), .D(
        OR4_1353_Y), .Y(OR4_348_Y));
    OR4 OR4_1098 (.A(\R_DATA_TEMPR80[21] ), .B(\R_DATA_TEMPR81[21] ), 
        .C(\R_DATA_TEMPR82[21] ), .D(\R_DATA_TEMPR83[21] ), .Y(
        OR4_1098_Y));
    OR4 OR4_162 (.A(\R_DATA_TEMPR120[28] ), .B(\R_DATA_TEMPR121[28] ), 
        .C(\R_DATA_TEMPR122[28] ), .D(\R_DATA_TEMPR123[28] ), .Y(
        OR4_162_Y));
    OR4 OR4_1387 (.A(OR4_1298_Y), .B(OR4_1102_Y), .C(OR4_734_Y), .D(
        OR4_578_Y), .Y(OR4_1387_Y));
    OR4 OR4_282 (.A(\R_DATA_TEMPR80[0] ), .B(\R_DATA_TEMPR81[0] ), .C(
        \R_DATA_TEMPR82[0] ), .D(\R_DATA_TEMPR83[0] ), .Y(OR4_282_Y));
    OR4 OR4_965 (.A(\R_DATA_TEMPR28[38] ), .B(\R_DATA_TEMPR29[38] ), 
        .C(\R_DATA_TEMPR30[38] ), .D(\R_DATA_TEMPR31[38] ), .Y(
        OR4_965_Y));
    OR4 OR4_316 (.A(\R_DATA_TEMPR76[28] ), .B(\R_DATA_TEMPR77[28] ), 
        .C(\R_DATA_TEMPR78[28] ), .D(\R_DATA_TEMPR79[28] ), .Y(
        OR4_316_Y));
    OR4 OR4_1612 (.A(\R_DATA_TEMPR40[21] ), .B(\R_DATA_TEMPR41[21] ), 
        .C(\R_DATA_TEMPR42[21] ), .D(\R_DATA_TEMPR43[21] ), .Y(
        OR4_1612_Y));
    OR4 OR4_1416 (.A(OR4_599_Y), .B(OR4_1624_Y), .C(OR4_236_Y), .D(
        OR4_805_Y), .Y(OR4_1416_Y));
    OR4 OR4_1314 (.A(\R_DATA_TEMPR24[12] ), .B(\R_DATA_TEMPR25[12] ), 
        .C(\R_DATA_TEMPR26[12] ), .D(\R_DATA_TEMPR27[12] ), .Y(
        OR4_1314_Y));
    OR4 OR4_909 (.A(\R_DATA_TEMPR88[17] ), .B(\R_DATA_TEMPR89[17] ), 
        .C(\R_DATA_TEMPR90[17] ), .D(\R_DATA_TEMPR91[17] ), .Y(
        OR4_909_Y));
    OR4 OR4_900 (.A(\R_DATA_TEMPR36[16] ), .B(\R_DATA_TEMPR37[16] ), 
        .C(\R_DATA_TEMPR38[16] ), .D(\R_DATA_TEMPR39[16] ), .Y(
        OR4_900_Y));
    OR4 OR4_1405 (.A(\R_DATA_TEMPR52[12] ), .B(\R_DATA_TEMPR53[12] ), 
        .C(\R_DATA_TEMPR54[12] ), .D(\R_DATA_TEMPR55[12] ), .Y(
        OR4_1405_Y));
    OR4 OR4_134 (.A(\R_DATA_TEMPR124[34] ), .B(\R_DATA_TEMPR125[34] ), 
        .C(\R_DATA_TEMPR126[34] ), .D(\R_DATA_TEMPR127[34] ), .Y(
        OR4_134_Y));
    OR4 OR4_1433 (.A(\R_DATA_TEMPR100[22] ), .B(\R_DATA_TEMPR101[22] ), 
        .C(\R_DATA_TEMPR102[22] ), .D(\R_DATA_TEMPR103[22] ), .Y(
        OR4_1433_Y));
    OR4 OR4_1592 (.A(\R_DATA_TEMPR68[11] ), .B(\R_DATA_TEMPR69[11] ), 
        .C(\R_DATA_TEMPR70[11] ), .D(\R_DATA_TEMPR71[11] ), .Y(
        OR4_1592_Y));
    OR4 OR4_723 (.A(\R_DATA_TEMPR56[8] ), .B(\R_DATA_TEMPR57[8] ), .C(
        \R_DATA_TEMPR58[8] ), .D(\R_DATA_TEMPR59[8] ), .Y(OR4_723_Y));
    OR2 OR2_35 (.A(\R_DATA_TEMPR84[26] ), .B(\R_DATA_TEMPR85[26] ), .Y(
        OR2_35_Y));
    OR4 OR4_979 (.A(OR4_1429_Y), .B(OR4_517_Y), .C(OR4_490_Y), .D(
        OR4_1263_Y), .Y(OR4_979_Y));
    OR4 OR4_970 (.A(\R_DATA_TEMPR92[28] ), .B(\R_DATA_TEMPR93[28] ), 
        .C(\R_DATA_TEMPR94[28] ), .D(\R_DATA_TEMPR95[28] ), .Y(
        OR4_970_Y));
    OR4 OR4_1067 (.A(\R_DATA_TEMPR108[25] ), .B(\R_DATA_TEMPR109[25] ), 
        .C(\R_DATA_TEMPR110[25] ), .D(\R_DATA_TEMPR111[25] ), .Y(
        OR4_1067_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%26%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C0 (.A_DOUT({
        \R_DATA_TEMPR26[39] , \R_DATA_TEMPR26[38] , 
        \R_DATA_TEMPR26[37] , \R_DATA_TEMPR26[36] , 
        \R_DATA_TEMPR26[35] , \R_DATA_TEMPR26[34] , 
        \R_DATA_TEMPR26[33] , \R_DATA_TEMPR26[32] , 
        \R_DATA_TEMPR26[31] , \R_DATA_TEMPR26[30] , 
        \R_DATA_TEMPR26[29] , \R_DATA_TEMPR26[28] , 
        \R_DATA_TEMPR26[27] , \R_DATA_TEMPR26[26] , 
        \R_DATA_TEMPR26[25] , \R_DATA_TEMPR26[24] , 
        \R_DATA_TEMPR26[23] , \R_DATA_TEMPR26[22] , 
        \R_DATA_TEMPR26[21] , \R_DATA_TEMPR26[20] }), .B_DOUT({
        \R_DATA_TEMPR26[19] , \R_DATA_TEMPR26[18] , 
        \R_DATA_TEMPR26[17] , \R_DATA_TEMPR26[16] , 
        \R_DATA_TEMPR26[15] , \R_DATA_TEMPR26[14] , 
        \R_DATA_TEMPR26[13] , \R_DATA_TEMPR26[12] , 
        \R_DATA_TEMPR26[11] , \R_DATA_TEMPR26[10] , 
        \R_DATA_TEMPR26[9] , \R_DATA_TEMPR26[8] , \R_DATA_TEMPR26[7] , 
        \R_DATA_TEMPR26[6] , \R_DATA_TEMPR26[5] , \R_DATA_TEMPR26[4] , 
        \R_DATA_TEMPR26[3] , \R_DATA_TEMPR26[2] , \R_DATA_TEMPR26[1] , 
        \R_DATA_TEMPR26[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_103 (.A(\R_DATA_TEMPR8[11] ), .B(\R_DATA_TEMPR9[11] ), .C(
        \R_DATA_TEMPR10[11] ), .D(\R_DATA_TEMPR11[11] ), .Y(OR4_103_Y));
    OR4 OR4_224 (.A(\R_DATA_TEMPR20[25] ), .B(\R_DATA_TEMPR21[25] ), 
        .C(\R_DATA_TEMPR22[25] ), .D(\R_DATA_TEMPR23[25] ), .Y(
        OR4_224_Y));
    OR4 OR4_149 (.A(\R_DATA_TEMPR36[15] ), .B(\R_DATA_TEMPR37[15] ), 
        .C(\R_DATA_TEMPR38[15] ), .D(\R_DATA_TEMPR39[15] ), .Y(
        OR4_149_Y));
    OR4 OR4_792 (.A(\R_DATA_TEMPR120[9] ), .B(\R_DATA_TEMPR121[9] ), 
        .C(\R_DATA_TEMPR122[9] ), .D(\R_DATA_TEMPR123[9] ), .Y(
        OR4_792_Y));
    OR4 OR4_380 (.A(\R_DATA_TEMPR92[38] ), .B(\R_DATA_TEMPR93[38] ), 
        .C(\R_DATA_TEMPR94[38] ), .D(\R_DATA_TEMPR95[38] ), .Y(
        OR4_380_Y));
    OR4 OR4_1617 (.A(\R_DATA_TEMPR36[30] ), .B(\R_DATA_TEMPR37[30] ), 
        .C(\R_DATA_TEMPR38[30] ), .D(\R_DATA_TEMPR39[30] ), .Y(
        OR4_1617_Y));
    OR4 OR4_933 (.A(\R_DATA_TEMPR64[24] ), .B(\R_DATA_TEMPR65[24] ), 
        .C(\R_DATA_TEMPR66[24] ), .D(\R_DATA_TEMPR67[24] ), .Y(
        OR4_933_Y));
    OR4 \OR4_R_DATA[13]  (.A(OR4_989_Y), .B(OR4_577_Y), .C(OR4_515_Y), 
        .D(OR4_465_Y), .Y(R_DATA[13]));
    OR4 OR4_173 (.A(\R_DATA_TEMPR16[30] ), .B(\R_DATA_TEMPR17[30] ), 
        .C(\R_DATA_TEMPR18[30] ), .D(\R_DATA_TEMPR19[30] ), .Y(
        OR4_173_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%33%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R33C0 (.A_DOUT({
        \R_DATA_TEMPR33[39] , \R_DATA_TEMPR33[38] , 
        \R_DATA_TEMPR33[37] , \R_DATA_TEMPR33[36] , 
        \R_DATA_TEMPR33[35] , \R_DATA_TEMPR33[34] , 
        \R_DATA_TEMPR33[33] , \R_DATA_TEMPR33[32] , 
        \R_DATA_TEMPR33[31] , \R_DATA_TEMPR33[30] , 
        \R_DATA_TEMPR33[29] , \R_DATA_TEMPR33[28] , 
        \R_DATA_TEMPR33[27] , \R_DATA_TEMPR33[26] , 
        \R_DATA_TEMPR33[25] , \R_DATA_TEMPR33[24] , 
        \R_DATA_TEMPR33[23] , \R_DATA_TEMPR33[22] , 
        \R_DATA_TEMPR33[21] , \R_DATA_TEMPR33[20] }), .B_DOUT({
        \R_DATA_TEMPR33[19] , \R_DATA_TEMPR33[18] , 
        \R_DATA_TEMPR33[17] , \R_DATA_TEMPR33[16] , 
        \R_DATA_TEMPR33[15] , \R_DATA_TEMPR33[14] , 
        \R_DATA_TEMPR33[13] , \R_DATA_TEMPR33[12] , 
        \R_DATA_TEMPR33[11] , \R_DATA_TEMPR33[10] , 
        \R_DATA_TEMPR33[9] , \R_DATA_TEMPR33[8] , \R_DATA_TEMPR33[7] , 
        \R_DATA_TEMPR33[6] , \R_DATA_TEMPR33[5] , \R_DATA_TEMPR33[4] , 
        \R_DATA_TEMPR33[3] , \R_DATA_TEMPR33[2] , \R_DATA_TEMPR33[1] , 
        \R_DATA_TEMPR33[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[33][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[8] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[8] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_269 (.A(OR4_741_Y), .B(OR4_1297_Y), .C(OR4_1155_Y), .D(
        OR4_499_Y), .Y(OR4_269_Y));
    OR4 OR4_996 (.A(\R_DATA_TEMPR100[26] ), .B(\R_DATA_TEMPR101[26] ), 
        .C(\R_DATA_TEMPR102[26] ), .D(\R_DATA_TEMPR103[26] ), .Y(
        OR4_996_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[31]  (.A(CFG3_23_Y), .B(
        CFG3_7_Y), .Y(\BLKX2[31] ));
    OR4 OR4_836 (.A(\R_DATA_TEMPR88[5] ), .B(\R_DATA_TEMPR89[5] ), .C(
        \R_DATA_TEMPR90[5] ), .D(\R_DATA_TEMPR91[5] ), .Y(OR4_836_Y));
    OR4 OR4_731 (.A(\R_DATA_TEMPR104[11] ), .B(\R_DATA_TEMPR105[11] ), 
        .C(\R_DATA_TEMPR106[11] ), .D(\R_DATA_TEMPR107[11] ), .Y(
        OR4_731_Y));
    OR4 OR4_695 (.A(\R_DATA_TEMPR24[33] ), .B(\R_DATA_TEMPR25[33] ), 
        .C(\R_DATA_TEMPR26[33] ), .D(\R_DATA_TEMPR27[33] ), .Y(
        OR4_695_Y));
    OR4 OR4_62 (.A(\R_DATA_TEMPR92[17] ), .B(\R_DATA_TEMPR93[17] ), .C(
        \R_DATA_TEMPR94[17] ), .D(\R_DATA_TEMPR95[17] ), .Y(OR4_62_Y));
    OR4 OR4_1604 (.A(\R_DATA_TEMPR16[25] ), .B(\R_DATA_TEMPR17[25] ), 
        .C(\R_DATA_TEMPR18[25] ), .D(\R_DATA_TEMPR19[25] ), .Y(
        OR4_1604_Y));
    OR4 OR4_883 (.A(\R_DATA_TEMPR108[17] ), .B(\R_DATA_TEMPR109[17] ), 
        .C(\R_DATA_TEMPR110[17] ), .D(\R_DATA_TEMPR111[17] ), .Y(
        OR4_883_Y));
    OR4 OR4_1175 (.A(\R_DATA_TEMPR76[36] ), .B(\R_DATA_TEMPR77[36] ), 
        .C(\R_DATA_TEMPR78[36] ), .D(\R_DATA_TEMPR79[36] ), .Y(
        OR4_1175_Y));
    OR4 OR4_941 (.A(OR4_653_Y), .B(OR4_151_Y), .C(OR4_126_Y), .D(
        OR4_1469_Y), .Y(OR4_941_Y));
    OR4 OR4_1485 (.A(\R_DATA_TEMPR68[1] ), .B(\R_DATA_TEMPR69[1] ), .C(
        \R_DATA_TEMPR70[1] ), .D(\R_DATA_TEMPR71[1] ), .Y(OR4_1485_Y));
    OR4 OR4_1319 (.A(\R_DATA_TEMPR8[12] ), .B(\R_DATA_TEMPR9[12] ), .C(
        \R_DATA_TEMPR10[12] ), .D(\R_DATA_TEMPR11[12] ), .Y(OR4_1319_Y)
        );
    OR4 OR4_38 (.A(OR4_355_Y), .B(OR4_82_Y), .C(OR4_1440_Y), .D(
        OR4_617_Y), .Y(OR4_38_Y));
    OR4 OR4_1250 (.A(OR4_172_Y), .B(OR4_1325_Y), .C(OR4_1373_Y), .D(
        OR4_573_Y), .Y(OR4_1250_Y));
    OR4 OR4_1071 (.A(OR4_1407_Y), .B(OR4_1152_Y), .C(OR4_70_Y), .D(
        OR4_526_Y), .Y(OR4_1071_Y));
    OR4 OR4_1010 (.A(\R_DATA_TEMPR32[38] ), .B(\R_DATA_TEMPR33[38] ), 
        .C(\R_DATA_TEMPR34[38] ), .D(\R_DATA_TEMPR35[38] ), .Y(
        OR4_1010_Y));
    OR4 OR4_325 (.A(\R_DATA_TEMPR68[16] ), .B(\R_DATA_TEMPR69[16] ), 
        .C(\R_DATA_TEMPR70[16] ), .D(\R_DATA_TEMPR71[16] ), .Y(
        OR4_325_Y));
    OR4 OR4_1306 (.A(\R_DATA_TEMPR20[26] ), .B(\R_DATA_TEMPR21[26] ), 
        .C(\R_DATA_TEMPR22[26] ), .D(\R_DATA_TEMPR23[26] ), .Y(
        OR4_1306_Y));
    OR4 OR4_536 (.A(\R_DATA_TEMPR44[10] ), .B(\R_DATA_TEMPR45[10] ), 
        .C(\R_DATA_TEMPR46[10] ), .D(\R_DATA_TEMPR47[10] ), .Y(
        OR4_536_Y));
    OR4 OR4_869 (.A(\R_DATA_TEMPR48[25] ), .B(\R_DATA_TEMPR49[25] ), 
        .C(\R_DATA_TEMPR50[25] ), .D(\R_DATA_TEMPR51[25] ), .Y(
        OR4_869_Y));
    OR4 OR4_1557 (.A(OR4_223_Y), .B(OR4_1176_Y), .C(OR4_1523_Y), .D(
        OR4_701_Y), .Y(OR4_1557_Y));
    OR4 OR4_1601 (.A(\R_DATA_TEMPR4[32] ), .B(\R_DATA_TEMPR5[32] ), .C(
        \R_DATA_TEMPR6[32] ), .D(\R_DATA_TEMPR7[32] ), .Y(OR4_1601_Y));
    OR4 OR4_1352 (.A(\R_DATA_TEMPR116[7] ), .B(\R_DATA_TEMPR117[7] ), 
        .C(\R_DATA_TEMPR118[7] ), .D(\R_DATA_TEMPR119[7] ), .Y(
        OR4_1352_Y));
    OR4 OR4_114 (.A(\R_DATA_TEMPR16[36] ), .B(\R_DATA_TEMPR17[36] ), 
        .C(\R_DATA_TEMPR18[36] ), .D(\R_DATA_TEMPR19[36] ), .Y(
        OR4_114_Y));
    OR4 OR4_155 (.A(\R_DATA_TEMPR60[23] ), .B(\R_DATA_TEMPR61[23] ), 
        .C(\R_DATA_TEMPR62[23] ), .D(\R_DATA_TEMPR63[23] ), .Y(
        OR4_155_Y));
    OR4 OR4_1423 (.A(\R_DATA_TEMPR92[3] ), .B(\R_DATA_TEMPR93[3] ), .C(
        \R_DATA_TEMPR94[3] ), .D(\R_DATA_TEMPR95[3] ), .Y(OR4_1423_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[6]  (.A(CFG3_10_Y), .B(
        CFG3_12_Y), .Y(\BLKX2[6] ));
    OR4 OR4_1252 (.A(OR4_192_Y), .B(OR4_497_Y), .C(OR4_203_Y), .D(
        OR4_1040_Y), .Y(OR4_1252_Y));
    OR4 OR4_800 (.A(OR4_1086_Y), .B(OR4_1352_Y), .C(OR4_1533_Y), .D(
        OR4_1526_Y), .Y(OR4_800_Y));
    OR4 OR4_1097 (.A(\R_DATA_TEMPR36[36] ), .B(\R_DATA_TEMPR37[36] ), 
        .C(\R_DATA_TEMPR38[36] ), .D(\R_DATA_TEMPR39[36] ), .Y(
        OR4_1097_Y));
    OR4 OR4_1073 (.A(\R_DATA_TEMPR48[12] ), .B(\R_DATA_TEMPR49[12] ), 
        .C(\R_DATA_TEMPR50[12] ), .D(\R_DATA_TEMPR51[12] ), .Y(
        OR4_1073_Y));
    OR4 OR4_1600 (.A(\R_DATA_TEMPR80[38] ), .B(\R_DATA_TEMPR81[38] ), 
        .C(\R_DATA_TEMPR82[38] ), .D(\R_DATA_TEMPR83[38] ), .Y(
        OR4_1600_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[14]  (.A(CFG3_10_Y), .B(
        CFG3_4_Y), .Y(\BLKX2[14] ));
    OR4 OR4_457 (.A(\R_DATA_TEMPR24[4] ), .B(\R_DATA_TEMPR25[4] ), .C(
        \R_DATA_TEMPR26[4] ), .D(\R_DATA_TEMPR27[4] ), .Y(OR4_457_Y));
    OR4 OR4_102 (.A(\R_DATA_TEMPR0[20] ), .B(\R_DATA_TEMPR1[20] ), .C(
        \R_DATA_TEMPR2[20] ), .D(\R_DATA_TEMPR3[20] ), .Y(OR4_102_Y));
    OR4 OR4_1419 (.A(\R_DATA_TEMPR76[18] ), .B(\R_DATA_TEMPR77[18] ), 
        .C(\R_DATA_TEMPR78[18] ), .D(\R_DATA_TEMPR79[18] ), .Y(
        OR4_1419_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[25]  (.A(CFG3_15_Y), .B(
        CFG3_3_Y), .Y(\BLKY2[25] ));
    OR4 OR4_1472 (.A(\R_DATA_TEMPR112[1] ), .B(\R_DATA_TEMPR113[1] ), 
        .C(\R_DATA_TEMPR114[1] ), .D(\R_DATA_TEMPR115[1] ), .Y(
        OR4_1472_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%107%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R107C0 (.A_DOUT({
        \R_DATA_TEMPR107[39] , \R_DATA_TEMPR107[38] , 
        \R_DATA_TEMPR107[37] , \R_DATA_TEMPR107[36] , 
        \R_DATA_TEMPR107[35] , \R_DATA_TEMPR107[34] , 
        \R_DATA_TEMPR107[33] , \R_DATA_TEMPR107[32] , 
        \R_DATA_TEMPR107[31] , \R_DATA_TEMPR107[30] , 
        \R_DATA_TEMPR107[29] , \R_DATA_TEMPR107[28] , 
        \R_DATA_TEMPR107[27] , \R_DATA_TEMPR107[26] , 
        \R_DATA_TEMPR107[25] , \R_DATA_TEMPR107[24] , 
        \R_DATA_TEMPR107[23] , \R_DATA_TEMPR107[22] , 
        \R_DATA_TEMPR107[21] , \R_DATA_TEMPR107[20] }), .B_DOUT({
        \R_DATA_TEMPR107[19] , \R_DATA_TEMPR107[18] , 
        \R_DATA_TEMPR107[17] , \R_DATA_TEMPR107[16] , 
        \R_DATA_TEMPR107[15] , \R_DATA_TEMPR107[14] , 
        \R_DATA_TEMPR107[13] , \R_DATA_TEMPR107[12] , 
        \R_DATA_TEMPR107[11] , \R_DATA_TEMPR107[10] , 
        \R_DATA_TEMPR107[9] , \R_DATA_TEMPR107[8] , 
        \R_DATA_TEMPR107[7] , \R_DATA_TEMPR107[6] , 
        \R_DATA_TEMPR107[5] , \R_DATA_TEMPR107[4] , 
        \R_DATA_TEMPR107[3] , \R_DATA_TEMPR107[2] , 
        \R_DATA_TEMPR107[1] , \R_DATA_TEMPR107[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[107][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[26] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[26] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_905 (.A(OR4_88_Y), .B(OR4_1546_Y), .C(OR4_43_Y), .D(
        OR4_654_Y), .Y(OR4_905_Y));
    OR4 OR4_870 (.A(\R_DATA_TEMPR24[20] ), .B(\R_DATA_TEMPR25[20] ), 
        .C(\R_DATA_TEMPR26[20] ), .D(\R_DATA_TEMPR27[20] ), .Y(
        OR4_870_Y));
    CFG1 #( .INIT(2'h1) )  \INVBLKY0[0]  (.A(R_ADDR[9]), .Y(\BLKY0[0] )
        );
    OR4 OR4_913 (.A(\R_DATA_TEMPR68[4] ), .B(\R_DATA_TEMPR69[4] ), .C(
        \R_DATA_TEMPR70[4] ), .D(\R_DATA_TEMPR71[4] ), .Y(OR4_913_Y));
    OR4 OR4_1454 (.A(\R_DATA_TEMPR60[30] ), .B(\R_DATA_TEMPR61[30] ), 
        .C(\R_DATA_TEMPR62[30] ), .D(\R_DATA_TEMPR63[30] ), .Y(
        OR4_1454_Y));
    OR4 OR4_690 (.A(\R_DATA_TEMPR88[34] ), .B(\R_DATA_TEMPR89[34] ), 
        .C(\R_DATA_TEMPR90[34] ), .D(\R_DATA_TEMPR91[34] ), .Y(
        OR4_690_Y));
    OR4 OR4_1133 (.A(\R_DATA_TEMPR56[0] ), .B(\R_DATA_TEMPR57[0] ), .C(
        \R_DATA_TEMPR58[0] ), .D(\R_DATA_TEMPR59[0] ), .Y(OR4_1133_Y));
    OR4 OR4_722 (.A(OR4_709_Y), .B(OR4_459_Y), .C(OR4_159_Y), .D(
        OR4_470_Y), .Y(OR4_722_Y));
    OR4 OR4_172 (.A(\R_DATA_TEMPR64[39] ), .B(\R_DATA_TEMPR65[39] ), 
        .C(\R_DATA_TEMPR66[39] ), .D(\R_DATA_TEMPR67[39] ), .Y(
        OR4_172_Y));
    OR4 OR4_745 (.A(\R_DATA_TEMPR64[21] ), .B(\R_DATA_TEMPR65[21] ), 
        .C(\R_DATA_TEMPR66[21] ), .D(\R_DATA_TEMPR67[21] ), .Y(
        OR4_745_Y));
    OR4 OR4_647 (.A(\R_DATA_TEMPR104[14] ), .B(\R_DATA_TEMPR105[14] ), 
        .C(\R_DATA_TEMPR106[14] ), .D(\R_DATA_TEMPR107[14] ), .Y(
        OR4_647_Y));
    OR4 OR4_1386 (.A(\R_DATA_TEMPR12[22] ), .B(\R_DATA_TEMPR13[22] ), 
        .C(\R_DATA_TEMPR14[22] ), .D(\R_DATA_TEMPR15[22] ), .Y(
        OR4_1386_Y));
    OR4 OR4_975 (.A(\R_DATA_TEMPR56[21] ), .B(\R_DATA_TEMPR57[21] ), 
        .C(\R_DATA_TEMPR58[21] ), .D(\R_DATA_TEMPR59[21] ), .Y(
        OR4_975_Y));
    OR4 OR4_1254 (.A(\R_DATA_TEMPR76[33] ), .B(\R_DATA_TEMPR77[33] ), 
        .C(\R_DATA_TEMPR78[33] ), .D(\R_DATA_TEMPR79[33] ), .Y(
        OR4_1254_Y));
    OR4 OR4_816 (.A(OR4_95_Y), .B(OR4_1559_Y), .C(OR4_53_Y), .D(
        OR4_312_Y), .Y(OR4_816_Y));
    OR4 OR4_746 (.A(\R_DATA_TEMPR76[4] ), .B(\R_DATA_TEMPR77[4] ), .C(
        \R_DATA_TEMPR78[4] ), .D(\R_DATA_TEMPR79[4] ), .Y(OR4_746_Y));
    OR4 OR4_711 (.A(\R_DATA_TEMPR92[1] ), .B(\R_DATA_TEMPR93[1] ), .C(
        \R_DATA_TEMPR94[1] ), .D(\R_DATA_TEMPR95[1] ), .Y(OR4_711_Y));
    OR4 OR4_585 (.A(\R_DATA_TEMPR68[29] ), .B(\R_DATA_TEMPR69[29] ), 
        .C(\R_DATA_TEMPR70[29] ), .D(\R_DATA_TEMPR71[29] ), .Y(
        OR4_585_Y));
    OR4 OR4_926 (.A(\R_DATA_TEMPR112[16] ), .B(\R_DATA_TEMPR113[16] ), 
        .C(\R_DATA_TEMPR114[16] ), .D(\R_DATA_TEMPR115[16] ), .Y(
        OR4_926_Y));
    OR4 OR4_767 (.A(OR4_703_Y), .B(OR4_447_Y), .C(OR4_148_Y), .D(
        OR4_1166_Y), .Y(OR4_767_Y));
    OR4 OR4_255 (.A(\R_DATA_TEMPR56[34] ), .B(\R_DATA_TEMPR57[34] ), 
        .C(\R_DATA_TEMPR58[34] ), .D(\R_DATA_TEMPR59[34] ), .Y(
        OR4_255_Y));
    OR4 OR4_397 (.A(OR4_773_Y), .B(OR4_1561_Y), .C(OR4_1535_Y), .D(
        OR4_1217_Y), .Y(OR4_397_Y));
    OR4 OR4_190 (.A(\R_DATA_TEMPR12[18] ), .B(\R_DATA_TEMPR13[18] ), 
        .C(\R_DATA_TEMPR14[18] ), .D(\R_DATA_TEMPR15[18] ), .Y(
        OR4_190_Y));
    OR4 OR4_1357 (.A(\R_DATA_TEMPR108[6] ), .B(\R_DATA_TEMPR109[6] ), 
        .C(\R_DATA_TEMPR110[6] ), .D(\R_DATA_TEMPR111[6] ), .Y(
        OR4_1357_Y));
    OR4 OR4_764 (.A(\R_DATA_TEMPR120[29] ), .B(\R_DATA_TEMPR121[29] ), 
        .C(\R_DATA_TEMPR122[29] ), .D(\R_DATA_TEMPR123[29] ), .Y(
        OR4_764_Y));
    OR4 OR4_1539 (.A(OR4_251_Y), .B(OR4_1399_Y), .C(OR4_294_Y), .D(
        OR4_739_Y), .Y(OR4_1539_Y));
    OR4 OR4_1408 (.A(\R_DATA_TEMPR44[19] ), .B(\R_DATA_TEMPR45[19] ), 
        .C(\R_DATA_TEMPR46[19] ), .D(\R_DATA_TEMPR47[19] ), .Y(
        OR4_1408_Y));
    OR4 OR4_625 (.A(OR4_1425_Y), .B(OR4_922_Y), .C(OR4_1006_Y), .D(
        OR4_1315_Y), .Y(OR4_625_Y));
    OR4 OR4_852 (.A(OR4_1074_Y), .B(OR4_1339_Y), .C(OR4_1522_Y), .D(
        OR4_1303_Y), .Y(OR4_852_Y));
    OR4 OR4_538 (.A(\R_DATA_TEMPR4[30] ), .B(\R_DATA_TEMPR5[30] ), .C(
        \R_DATA_TEMPR6[30] ), .D(\R_DATA_TEMPR7[30] ), .Y(OR4_538_Y));
    OR4 OR4_26 (.A(\R_DATA_TEMPR100[25] ), .B(\R_DATA_TEMPR101[25] ), 
        .C(\R_DATA_TEMPR102[25] ), .D(\R_DATA_TEMPR103[25] ), .Y(
        OR4_26_Y));
    OR4 OR4_53 (.A(\R_DATA_TEMPR120[18] ), .B(\R_DATA_TEMPR121[18] ), 
        .C(\R_DATA_TEMPR122[18] ), .D(\R_DATA_TEMPR123[18] ), .Y(
        OR4_53_Y));
    OR4 OR4_683 (.A(\R_DATA_TEMPR112[19] ), .B(\R_DATA_TEMPR113[19] ), 
        .C(\R_DATA_TEMPR114[19] ), .D(\R_DATA_TEMPR115[19] ), .Y(
        OR4_683_Y));
    OR4 OR4_209 (.A(\R_DATA_TEMPR4[2] ), .B(\R_DATA_TEMPR5[2] ), .C(
        \R_DATA_TEMPR6[2] ), .D(\R_DATA_TEMPR7[2] ), .Y(OR4_209_Y));
    OR4 OR4_798 (.A(OR4_220_Y), .B(OR2_39_Y), .C(\R_DATA_TEMPR86[31] ), 
        .D(\R_DATA_TEMPR87[31] ), .Y(OR4_798_Y));
    OR4 OR4_861 (.A(OR4_93_Y), .B(OR4_1555_Y), .C(OR4_48_Y), .D(
        OR4_1575_Y), .Y(OR4_861_Y));
    OR4 OR4_516 (.A(OR4_869_Y), .B(OR4_1459_Y), .C(OR4_601_Y), .D(
        OR4_859_Y), .Y(OR4_516_Y));
    OR4 OR4_279 (.A(\R_DATA_TEMPR52[35] ), .B(\R_DATA_TEMPR53[35] ), 
        .C(\R_DATA_TEMPR54[35] ), .D(\R_DATA_TEMPR55[35] ), .Y(
        OR4_279_Y));
    OR4 OR4_1267 (.A(\R_DATA_TEMPR72[31] ), .B(\R_DATA_TEMPR73[31] ), 
        .C(\R_DATA_TEMPR74[31] ), .D(\R_DATA_TEMPR75[31] ), .Y(
        OR4_1267_Y));
    OR4 OR4_436 (.A(OR4_1122_Y), .B(OR4_286_Y), .C(OR4_743_Y), .D(
        OR4_1048_Y), .Y(OR4_436_Y));
    OR4 OR4_89 (.A(\R_DATA_TEMPR108[12] ), .B(\R_DATA_TEMPR109[12] ), 
        .C(\R_DATA_TEMPR110[12] ), .D(\R_DATA_TEMPR111[12] ), .Y(
        OR4_89_Y));
    OR4 OR4_453 (.A(\R_DATA_TEMPR104[37] ), .B(\R_DATA_TEMPR105[37] ), 
        .C(\R_DATA_TEMPR106[37] ), .D(\R_DATA_TEMPR107[37] ), .Y(
        OR4_453_Y));
    OR4 OR4_1104 (.A(\R_DATA_TEMPR72[4] ), .B(\R_DATA_TEMPR73[4] ), .C(
        \R_DATA_TEMPR74[4] ), .D(\R_DATA_TEMPR75[4] ), .Y(OR4_1104_Y));
    OR4 OR4_897 (.A(\R_DATA_TEMPR92[12] ), .B(\R_DATA_TEMPR93[12] ), 
        .C(\R_DATA_TEMPR94[12] ), .D(\R_DATA_TEMPR95[12] ), .Y(
        OR4_897_Y));
    OR4 OR4_651 (.A(\R_DATA_TEMPR108[23] ), .B(\R_DATA_TEMPR109[23] ), 
        .C(\R_DATA_TEMPR110[23] ), .D(\R_DATA_TEMPR111[23] ), .Y(
        OR4_651_Y));
    OR4 OR4_198 (.A(\R_DATA_TEMPR80[22] ), .B(\R_DATA_TEMPR81[22] ), 
        .C(\R_DATA_TEMPR82[22] ), .D(\R_DATA_TEMPR83[22] ), .Y(
        OR4_198_Y));
    OR4 OR4_1410 (.A(\R_DATA_TEMPR120[8] ), .B(\R_DATA_TEMPR121[8] ), 
        .C(\R_DATA_TEMPR122[8] ), .D(\R_DATA_TEMPR123[8] ), .Y(
        OR4_1410_Y));
    OR4 OR4_1078 (.A(OR4_171_Y), .B(OR4_6_Y), .C(OR4_125_Y), .D(
        OR4_525_Y), .Y(OR4_1078_Y));
    OR4 OR4_994 (.A(\R_DATA_TEMPR8[28] ), .B(\R_DATA_TEMPR9[28] ), .C(
        \R_DATA_TEMPR10[28] ), .D(\R_DATA_TEMPR11[28] ), .Y(OR4_994_Y));
    OR4 OR4_1488 (.A(OR4_831_Y), .B(OR4_659_Y), .C(OR4_61_Y), .D(
        OR4_582_Y), .Y(OR4_1488_Y));
    OR4 OR4_989 (.A(OR4_1537_Y), .B(OR4_1211_Y), .C(OR4_1180_Y), .D(
        OR4_563_Y), .Y(OR4_989_Y));
    OR4 OR4_980 (.A(\R_DATA_TEMPR64[10] ), .B(\R_DATA_TEMPR65[10] ), 
        .C(\R_DATA_TEMPR66[10] ), .D(\R_DATA_TEMPR67[10] ), .Y(
        OR4_980_Y));
    OR4 OR4_809 (.A(OR4_1089_Y), .B(OR4_921_Y), .C(OR4_1477_Y), .D(
        OR4_292_Y), .Y(OR4_809_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[3]  (.A(CFG3_5_Y), .B(CFG3_12_Y)
        , .Y(\BLKX2[3] ));
    OR4 OR4_1544 (.A(OR4_528_Y), .B(OR4_826_Y), .C(OR4_1065_Y), .D(
        OR4_883_Y), .Y(OR4_1544_Y));
    OR4 OR4_258 (.A(\R_DATA_TEMPR120[21] ), .B(\R_DATA_TEMPR121[21] ), 
        .C(\R_DATA_TEMPR122[21] ), .D(\R_DATA_TEMPR123[21] ), .Y(
        OR4_258_Y));
    OR4 OR4_1466 (.A(OR4_1312_Y), .B(OR4_253_Y), .C(OR4_1024_Y), .D(
        OR4_1294_Y), .Y(OR4_1466_Y));
    OR4 OR4_1364 (.A(\R_DATA_TEMPR20[20] ), .B(\R_DATA_TEMPR21[20] ), 
        .C(\R_DATA_TEMPR22[20] ), .D(\R_DATA_TEMPR23[20] ), .Y(
        OR4_1364_Y));
    OR4 \OR4_R_DATA[21]  (.A(OR4_1505_Y), .B(OR4_1434_Y), .C(
        OR4_1466_Y), .D(OR4_937_Y), .Y(R_DATA[21]));
    OR4 OR4_1123 (.A(\R_DATA_TEMPR0[13] ), .B(\R_DATA_TEMPR1[13] ), .C(
        \R_DATA_TEMPR2[13] ), .D(\R_DATA_TEMPR3[13] ), .Y(OR4_1123_Y));
    OR4 OR4_1500 (.A(\R_DATA_TEMPR60[4] ), .B(\R_DATA_TEMPR61[4] ), .C(
        \R_DATA_TEMPR62[4] ), .D(\R_DATA_TEMPR63[4] ), .Y(OR4_1500_Y));
    OR4 OR4_1455 (.A(OR4_114_Y), .B(OR4_638_Y), .C(OR4_131_Y), .D(
        OR4_1276_Y), .Y(OR4_1455_Y));
    OR4 OR4_620 (.A(\R_DATA_TEMPR52[37] ), .B(\R_DATA_TEMPR53[37] ), 
        .C(\R_DATA_TEMPR54[37] ), .D(\R_DATA_TEMPR55[37] ), .Y(
        OR4_620_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[27]  (.A(CFG3_5_Y), .B(CFG3_7_Y)
        , .Y(\BLKX2[27] ));
    OR4 OR4_1345 (.A(\R_DATA_TEMPR4[4] ), .B(\R_DATA_TEMPR5[4] ), .C(
        \R_DATA_TEMPR6[4] ), .D(\R_DATA_TEMPR7[4] ), .Y(OR4_1345_Y));
    OR4 OR4_879 (.A(\R_DATA_TEMPR76[3] ), .B(\R_DATA_TEMPR77[3] ), .C(
        \R_DATA_TEMPR78[3] ), .D(\R_DATA_TEMPR79[3] ), .Y(OR4_879_Y));
    OR4 OR4_183 (.A(\R_DATA_TEMPR24[16] ), .B(\R_DATA_TEMPR25[16] ), 
        .C(\R_DATA_TEMPR26[16] ), .D(\R_DATA_TEMPR27[16] ), .Y(
        OR4_183_Y));
    OR4 OR4_1111 (.A(OR4_1547_Y), .B(OR4_1047_Y), .C(OR4_1105_Y), .D(
        OR4_1375_Y), .Y(OR4_1111_Y));
    OR4 OR4_332 (.A(OR4_980_Y), .B(OR4_817_Y), .C(OR4_938_Y), .D(
        OR4_777_Y), .Y(OR4_332_Y));
    OR4 OR4_1572 (.A(\R_DATA_TEMPR40[27] ), .B(\R_DATA_TEMPR41[27] ), 
        .C(\R_DATA_TEMPR42[27] ), .D(\R_DATA_TEMPR43[27] ), .Y(
        OR4_1572_Y));
    OR4 OR4_13 (.A(\R_DATA_TEMPR56[37] ), .B(\R_DATA_TEMPR57[37] ), .C(
        \R_DATA_TEMPR58[37] ), .D(\R_DATA_TEMPR59[37] ), .Y(OR4_13_Y));
    OR4 OR4_247 (.A(OR4_1390_Y), .B(OR4_1020_Y), .C(OR4_1572_Y), .D(
        OR4_959_Y), .Y(OR4_247_Y));
    OR4 OR4_1208 (.A(OR4_22_Y), .B(OR4_557_Y), .C(OR4_54_Y), .D(
        OR4_1181_Y), .Y(OR4_1208_Y));
    OR4 OR4_1529 (.A(OR4_971_Y), .B(OR4_1365_Y), .C(OR4_268_Y), .D(
        OR4_711_Y), .Y(OR4_1529_Y));
    CFG3 #( .INIT(8'h80) )  CFG3_3 (.A(R_EN), .B(R_ADDR[15]), .C(
        R_ADDR[14]), .Y(CFG3_3_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%125%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R125C0 (.A_DOUT({
        \R_DATA_TEMPR125[39] , \R_DATA_TEMPR125[38] , 
        \R_DATA_TEMPR125[37] , \R_DATA_TEMPR125[36] , 
        \R_DATA_TEMPR125[35] , \R_DATA_TEMPR125[34] , 
        \R_DATA_TEMPR125[33] , \R_DATA_TEMPR125[32] , 
        \R_DATA_TEMPR125[31] , \R_DATA_TEMPR125[30] , 
        \R_DATA_TEMPR125[29] , \R_DATA_TEMPR125[28] , 
        \R_DATA_TEMPR125[27] , \R_DATA_TEMPR125[26] , 
        \R_DATA_TEMPR125[25] , \R_DATA_TEMPR125[24] , 
        \R_DATA_TEMPR125[23] , \R_DATA_TEMPR125[22] , 
        \R_DATA_TEMPR125[21] , \R_DATA_TEMPR125[20] }), .B_DOUT({
        \R_DATA_TEMPR125[19] , \R_DATA_TEMPR125[18] , 
        \R_DATA_TEMPR125[17] , \R_DATA_TEMPR125[16] , 
        \R_DATA_TEMPR125[15] , \R_DATA_TEMPR125[14] , 
        \R_DATA_TEMPR125[13] , \R_DATA_TEMPR125[12] , 
        \R_DATA_TEMPR125[11] , \R_DATA_TEMPR125[10] , 
        \R_DATA_TEMPR125[9] , \R_DATA_TEMPR125[8] , 
        \R_DATA_TEMPR125[7] , \R_DATA_TEMPR125[6] , 
        \R_DATA_TEMPR125[5] , \R_DATA_TEMPR125[4] , 
        \R_DATA_TEMPR125[3] , \R_DATA_TEMPR125[2] , 
        \R_DATA_TEMPR125[1] , \R_DATA_TEMPR125[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[125][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[31] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[31] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_518 (.A(\R_DATA_TEMPR68[13] ), .B(\R_DATA_TEMPR69[13] ), 
        .C(\R_DATA_TEMPR70[13] ), .D(\R_DATA_TEMPR71[13] ), .Y(
        OR4_518_Y));
    OR4 OR4_147 (.A(\R_DATA_TEMPR52[2] ), .B(\R_DATA_TEMPR53[2] ), .C(
        \R_DATA_TEMPR54[2] ), .D(\R_DATA_TEMPR55[2] ), .Y(OR4_147_Y));
    OR4 OR4_327 (.A(\R_DATA_TEMPR28[5] ), .B(\R_DATA_TEMPR29[5] ), .C(
        \R_DATA_TEMPR30[5] ), .D(\R_DATA_TEMPR31[5] ), .Y(OR4_327_Y));
    OR4 OR4_120 (.A(\R_DATA_TEMPR48[11] ), .B(\R_DATA_TEMPR49[11] ), 
        .C(\R_DATA_TEMPR50[11] ), .D(\R_DATA_TEMPR51[11] ), .Y(
        OR4_120_Y));
    OR4 OR4_1535 (.A(\R_DATA_TEMPR88[36] ), .B(\R_DATA_TEMPR89[36] ), 
        .C(\R_DATA_TEMPR90[36] ), .D(\R_DATA_TEMPR91[36] ), .Y(
        OR4_1535_Y));
    OR4 OR4_1516 (.A(\R_DATA_TEMPR80[35] ), .B(\R_DATA_TEMPR81[35] ), 
        .C(\R_DATA_TEMPR82[35] ), .D(\R_DATA_TEMPR83[35] ), .Y(
        OR4_1516_Y));
    CFG1 #( .INIT(2'h1) )  \INVBLKY1[0]  (.A(R_ADDR[10]), .Y(
        \BLKY1[0] ));
    OR4 OR4_51 (.A(\R_DATA_TEMPR124[23] ), .B(\R_DATA_TEMPR125[23] ), 
        .C(\R_DATA_TEMPR126[23] ), .D(\R_DATA_TEMPR127[23] ), .Y(
        OR4_51_Y));
    OR4 OR4_967 (.A(\R_DATA_TEMPR120[3] ), .B(\R_DATA_TEMPR121[3] ), 
        .C(\R_DATA_TEMPR122[3] ), .D(\R_DATA_TEMPR123[3] ), .Y(
        OR4_967_Y));
    OR2 OR2_2 (.A(\R_DATA_TEMPR84[25] ), .B(\R_DATA_TEMPR85[25] ), .Y(
        OR2_2_Y));
    OR4 \OR4_R_DATA[20]  (.A(OR4_1195_Y), .B(OR4_1574_Y), .C(OR4_675_Y)
        , .D(OR4_55_Y), .Y(R_DATA[20]));
    OR4 OR4_1184 (.A(\R_DATA_TEMPR124[20] ), .B(\R_DATA_TEMPR125[20] ), 
        .C(\R_DATA_TEMPR126[20] ), .D(\R_DATA_TEMPR127[20] ), .Y(
        OR4_1184_Y));
    OR4 OR4_1236 (.A(OR4_1460_Y), .B(OR4_392_Y), .C(OR4_1161_Y), .D(
        OR4_1442_Y), .Y(OR4_1236_Y));
    OR4 OR4_728 (.A(\R_DATA_TEMPR40[31] ), .B(\R_DATA_TEMPR41[31] ), 
        .C(\R_DATA_TEMPR42[31] ), .D(\R_DATA_TEMPR43[31] ), .Y(
        OR4_728_Y));
    OR4 OR4_707 (.A(OR4_1395_Y), .B(OR4_3_Y), .C(OR4_200_Y), .D(
        OR4_367_Y), .Y(OR4_707_Y));
    OR4 OR4_1297 (.A(OR4_36_Y), .B(OR4_895_Y), .C(OR4_59_Y), .D(
        OR4_327_Y), .Y(OR4_1297_Y));
    OR4 OR4_704 (.A(\R_DATA_TEMPR40[14] ), .B(\R_DATA_TEMPR41[14] ), 
        .C(\R_DATA_TEMPR42[14] ), .D(\R_DATA_TEMPR43[14] ), .Y(
        OR4_704_Y));
    OR4 OR4_1580 (.A(\R_DATA_TEMPR88[28] ), .B(\R_DATA_TEMPR89[28] ), 
        .C(\R_DATA_TEMPR90[28] ), .D(\R_DATA_TEMPR91[28] ), .Y(
        OR4_1580_Y));
    OR4 OR4_1369 (.A(\R_DATA_TEMPR0[28] ), .B(\R_DATA_TEMPR1[28] ), .C(
        \R_DATA_TEMPR2[28] ), .D(\R_DATA_TEMPR3[28] ), .Y(OR4_1369_Y));
    OR2 OR2_39 (.A(\R_DATA_TEMPR84[31] ), .B(\R_DATA_TEMPR85[31] ), .Y(
        OR2_39_Y));
    OR4 OR4_20 (.A(OR4_733_Y), .B(OR4_1637_Y), .C(OR4_546_Y), .D(
        OR4_1571_Y), .Y(OR4_20_Y));
    OR4 OR4_1338 (.A(\R_DATA_TEMPR60[29] ), .B(\R_DATA_TEMPR61[29] ), 
        .C(\R_DATA_TEMPR62[29] ), .D(\R_DATA_TEMPR63[29] ), .Y(
        OR4_1338_Y));
    OR4 OR4_743 (.A(\R_DATA_TEMPR8[15] ), .B(\R_DATA_TEMPR9[15] ), .C(
        \R_DATA_TEMPR10[15] ), .D(\R_DATA_TEMPR11[15] ), .Y(OR4_743_Y));
    OR4 OR4_1060 (.A(\R_DATA_TEMPR36[21] ), .B(\R_DATA_TEMPR37[21] ), 
        .C(\R_DATA_TEMPR38[21] ), .D(\R_DATA_TEMPR39[21] ), .Y(
        OR4_1060_Y));
    OR4 OR4_777 (.A(\R_DATA_TEMPR76[10] ), .B(\R_DATA_TEMPR77[10] ), 
        .C(\R_DATA_TEMPR78[10] ), .D(\R_DATA_TEMPR79[10] ), .Y(
        OR4_777_Y));
    OR4 OR4_416 (.A(\R_DATA_TEMPR100[30] ), .B(\R_DATA_TEMPR101[30] ), 
        .C(\R_DATA_TEMPR102[30] ), .D(\R_DATA_TEMPR103[30] ), .Y(
        OR4_416_Y));
    OR4 \OR4_R_DATA[26]  (.A(OR4_625_Y), .B(OR4_1514_Y), .C(OR4_163_Y), 
        .D(OR4_261_Y), .Y(R_DATA[26]));
    OR4 OR4_774 (.A(\R_DATA_TEMPR60[34] ), .B(\R_DATA_TEMPR61[34] ), 
        .C(\R_DATA_TEMPR62[34] ), .D(\R_DATA_TEMPR63[34] ), .Y(
        OR4_774_Y));
    OR4 OR4_1417 (.A(\R_DATA_TEMPR92[6] ), .B(\R_DATA_TEMPR93[6] ), .C(
        \R_DATA_TEMPR94[6] ), .D(\R_DATA_TEMPR95[6] ), .Y(OR4_1417_Y));
    OR4 OR4_244 (.A(\R_DATA_TEMPR60[28] ), .B(\R_DATA_TEMPR61[28] ), 
        .C(\R_DATA_TEMPR62[28] ), .D(\R_DATA_TEMPR63[28] ), .Y(
        OR4_244_Y));
    OR4 OR4_1356 (.A(\R_DATA_TEMPR92[11] ), .B(\R_DATA_TEMPR93[11] ), 
        .C(\R_DATA_TEMPR94[11] ), .D(\R_DATA_TEMPR95[11] ), .Y(
        OR4_1356_Y));
    OR4 OR4_801 (.A(\R_DATA_TEMPR8[31] ), .B(\R_DATA_TEMPR9[31] ), .C(
        \R_DATA_TEMPR10[31] ), .D(\R_DATA_TEMPR11[31] ), .Y(OR4_801_Y));
    OR4 OR4_1288 (.A(OR4_311_Y), .B(OR4_1243_Y), .C(OR4_1323_Y), .D(
        OR4_516_Y), .Y(OR4_1288_Y));
    OR4 OR4_27 (.A(\R_DATA_TEMPR88[21] ), .B(\R_DATA_TEMPR89[21] ), .C(
        \R_DATA_TEMPR90[21] ), .D(\R_DATA_TEMPR91[21] ), .Y(OR4_27_Y));
    OR4 OR4_1496 (.A(\R_DATA_TEMPR104[16] ), .B(\R_DATA_TEMPR105[16] ), 
        .C(\R_DATA_TEMPR106[16] ), .D(\R_DATA_TEMPR107[16] ), .Y(
        OR4_1496_Y));
    OR4 OR4_1394 (.A(\R_DATA_TEMPR64[28] ), .B(\R_DATA_TEMPR65[28] ), 
        .C(\R_DATA_TEMPR66[28] ), .D(\R_DATA_TEMPR67[28] ), .Y(
        OR4_1394_Y));
    OR4 OR4_82 (.A(\R_DATA_TEMPR116[22] ), .B(\R_DATA_TEMPR117[22] ), 
        .C(\R_DATA_TEMPR118[22] ), .D(\R_DATA_TEMPR119[22] ), .Y(
        OR4_82_Y));
    OR4 OR4_827 (.A(OR4_1118_Y), .B(OR4_627_Y), .C(OR4_677_Y), .D(
        OR4_1376_Y), .Y(OR4_827_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%66%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R66C0 (.A_DOUT({
        \R_DATA_TEMPR66[39] , \R_DATA_TEMPR66[38] , 
        \R_DATA_TEMPR66[37] , \R_DATA_TEMPR66[36] , 
        \R_DATA_TEMPR66[35] , \R_DATA_TEMPR66[34] , 
        \R_DATA_TEMPR66[33] , \R_DATA_TEMPR66[32] , 
        \R_DATA_TEMPR66[31] , \R_DATA_TEMPR66[30] , 
        \R_DATA_TEMPR66[29] , \R_DATA_TEMPR66[28] , 
        \R_DATA_TEMPR66[27] , \R_DATA_TEMPR66[26] , 
        \R_DATA_TEMPR66[25] , \R_DATA_TEMPR66[24] , 
        \R_DATA_TEMPR66[23] , \R_DATA_TEMPR66[22] , 
        \R_DATA_TEMPR66[21] , \R_DATA_TEMPR66[20] }), .B_DOUT({
        \R_DATA_TEMPR66[19] , \R_DATA_TEMPR66[18] , 
        \R_DATA_TEMPR66[17] , \R_DATA_TEMPR66[16] , 
        \R_DATA_TEMPR66[15] , \R_DATA_TEMPR66[14] , 
        \R_DATA_TEMPR66[13] , \R_DATA_TEMPR66[12] , 
        \R_DATA_TEMPR66[11] , \R_DATA_TEMPR66[10] , 
        \R_DATA_TEMPR66[9] , \R_DATA_TEMPR66[8] , \R_DATA_TEMPR66[7] , 
        \R_DATA_TEMPR66[6] , \R_DATA_TEMPR66[5] , \R_DATA_TEMPR66[4] , 
        \R_DATA_TEMPR66[3] , \R_DATA_TEMPR66[2] , \R_DATA_TEMPR66[1] , 
        \R_DATA_TEMPR66[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[66][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[16] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[16] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_128 (.A(\R_DATA_TEMPR68[33] ), .B(\R_DATA_TEMPR69[33] ), 
        .C(\R_DATA_TEMPR70[33] ), .D(\R_DATA_TEMPR71[33] ), .Y(
        OR4_128_Y));
    OR4 OR4_230 (.A(\R_DATA_TEMPR92[19] ), .B(\R_DATA_TEMPR93[19] ), 
        .C(\R_DATA_TEMPR94[19] ), .D(\R_DATA_TEMPR95[19] ), .Y(
        OR4_230_Y));
    OR4 OR4_924 (.A(\R_DATA_TEMPR48[39] ), .B(\R_DATA_TEMPR49[39] ), 
        .C(\R_DATA_TEMPR50[39] ), .D(\R_DATA_TEMPR51[39] ), .Y(
        OR4_924_Y));
    OR4 OR4_1015 (.A(\R_DATA_TEMPR112[2] ), .B(\R_DATA_TEMPR113[2] ), 
        .C(\R_DATA_TEMPR114[2] ), .D(\R_DATA_TEMPR115[2] ), .Y(
        OR4_1015_Y));
    OR4 OR4_537 (.A(\R_DATA_TEMPR16[27] ), .B(\R_DATA_TEMPR17[27] ), 
        .C(\R_DATA_TEMPR18[27] ), .D(\R_DATA_TEMPR19[27] ), .Y(
        OR4_537_Y));
    OR4 OR4_880 (.A(\R_DATA_TEMPR20[0] ), .B(\R_DATA_TEMPR21[0] ), .C(
        \R_DATA_TEMPR22[0] ), .D(\R_DATA_TEMPR23[0] ), .Y(OR4_880_Y));
    OR4 OR4_871 (.A(\R_DATA_TEMPR40[16] ), .B(\R_DATA_TEMPR41[16] ), 
        .C(\R_DATA_TEMPR42[16] ), .D(\R_DATA_TEMPR43[16] ), .Y(
        OR4_871_Y));
    OR4 OR4_182 (.A(OR4_1610_Y), .B(OR4_1350_Y), .C(OR4_1055_Y), .D(
        OR4_1313_Y), .Y(OR4_182_Y));
    OR4 OR4_312 (.A(\R_DATA_TEMPR124[18] ), .B(\R_DATA_TEMPR125[18] ), 
        .C(\R_DATA_TEMPR126[18] ), .D(\R_DATA_TEMPR127[18] ), .Y(
        OR4_312_Y));
    OR4 OR4_465 (.A(OR4_1158_Y), .B(OR4_992_Y), .C(OR4_1120_Y), .D(
        OR4_1150_Y), .Y(OR4_465_Y));
    OR4 OR4_551 (.A(\R_DATA_TEMPR52[26] ), .B(\R_DATA_TEMPR53[26] ), 
        .C(\R_DATA_TEMPR54[26] ), .D(\R_DATA_TEMPR55[26] ), .Y(
        OR4_551_Y));
    OR4 OR4_64 (.A(\R_DATA_TEMPR52[0] ), .B(\R_DATA_TEMPR53[0] ), .C(
        \R_DATA_TEMPR54[0] ), .D(\R_DATA_TEMPR55[0] ), .Y(OR4_64_Y));
    OR4 OR4_1469 (.A(\R_DATA_TEMPR92[33] ), .B(\R_DATA_TEMPR93[33] ), 
        .C(\R_DATA_TEMPR94[33] ), .D(\R_DATA_TEMPR95[33] ), .Y(
        OR4_1469_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%74%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R74C0 (.A_DOUT({
        \R_DATA_TEMPR74[39] , \R_DATA_TEMPR74[38] , 
        \R_DATA_TEMPR74[37] , \R_DATA_TEMPR74[36] , 
        \R_DATA_TEMPR74[35] , \R_DATA_TEMPR74[34] , 
        \R_DATA_TEMPR74[33] , \R_DATA_TEMPR74[32] , 
        \R_DATA_TEMPR74[31] , \R_DATA_TEMPR74[30] , 
        \R_DATA_TEMPR74[29] , \R_DATA_TEMPR74[28] , 
        \R_DATA_TEMPR74[27] , \R_DATA_TEMPR74[26] , 
        \R_DATA_TEMPR74[25] , \R_DATA_TEMPR74[24] , 
        \R_DATA_TEMPR74[23] , \R_DATA_TEMPR74[22] , 
        \R_DATA_TEMPR74[21] , \R_DATA_TEMPR74[20] }), .B_DOUT({
        \R_DATA_TEMPR74[19] , \R_DATA_TEMPR74[18] , 
        \R_DATA_TEMPR74[17] , \R_DATA_TEMPR74[16] , 
        \R_DATA_TEMPR74[15] , \R_DATA_TEMPR74[14] , 
        \R_DATA_TEMPR74[13] , \R_DATA_TEMPR74[12] , 
        \R_DATA_TEMPR74[11] , \R_DATA_TEMPR74[10] , 
        \R_DATA_TEMPR74[9] , \R_DATA_TEMPR74[8] , \R_DATA_TEMPR74[7] , 
        \R_DATA_TEMPR74[6] , \R_DATA_TEMPR74[5] , \R_DATA_TEMPR74[4] , 
        \R_DATA_TEMPR74[3] , \R_DATA_TEMPR74[2] , \R_DATA_TEMPR74[1] , 
        \R_DATA_TEMPR74[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[74][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[18] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[18] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1609 (.A(\R_DATA_TEMPR20[34] ), .B(\R_DATA_TEMPR21[34] ), 
        .C(\R_DATA_TEMPR22[34] ), .D(\R_DATA_TEMPR23[34] ), .Y(
        OR4_1609_Y));
    OR4 OR4_1105 (.A(\R_DATA_TEMPR120[35] ), .B(\R_DATA_TEMPR121[35] ), 
        .C(\R_DATA_TEMPR122[35] ), .D(\R_DATA_TEMPR123[35] ), .Y(
        OR4_1105_Y));
    OR4 OR4_1077 (.A(OR4_45_Y), .B(OR4_368_Y), .C(OR4_1451_Y), .D(
        OR4_660_Y), .Y(OR4_1077_Y));
    OR4 OR4_985 (.A(\R_DATA_TEMPR20[28] ), .B(\R_DATA_TEMPR21[28] ), 
        .C(\R_DATA_TEMPR22[28] ), .D(\R_DATA_TEMPR23[28] ), .Y(
        OR4_985_Y));
    OR4 OR4_11 (.A(\R_DATA_TEMPR40[1] ), .B(\R_DATA_TEMPR41[1] ), .C(
        \R_DATA_TEMPR42[1] ), .D(\R_DATA_TEMPR43[1] ), .Y(OR4_11_Y));
    OR4 OR4_1039 (.A(\R_DATA_TEMPR76[13] ), .B(\R_DATA_TEMPR77[13] ), 
        .C(\R_DATA_TEMPR78[13] ), .D(\R_DATA_TEMPR79[13] ), .Y(
        OR4_1039_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[10]  (.A(CFG3_14_Y), .B(
        CFG3_4_Y), .Y(\BLKX2[10] ));
    OR4 OR4_639 (.A(\R_DATA_TEMPR72[13] ), .B(\R_DATA_TEMPR73[13] ), 
        .C(\R_DATA_TEMPR74[13] ), .D(\R_DATA_TEMPR75[13] ), .Y(
        OR4_639_Y));
    OR4 OR4_1001 (.A(\R_DATA_TEMPR56[32] ), .B(\R_DATA_TEMPR57[32] ), 
        .C(\R_DATA_TEMPR58[32] ), .D(\R_DATA_TEMPR59[32] ), .Y(
        OR4_1001_Y));
    OR4 OR4_1525 (.A(\R_DATA_TEMPR104[35] ), .B(\R_DATA_TEMPR105[35] ), 
        .C(\R_DATA_TEMPR106[35] ), .D(\R_DATA_TEMPR107[35] ), .Y(
        OR4_1525_Y));
    OR4 OR4_345 (.A(OR4_1073_Y), .B(OR4_1405_Y), .C(OR4_1636_Y), .D(
        OR4_1453_Y), .Y(OR4_345_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%84%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R84C0 (.A_DOUT({
        \R_DATA_TEMPR84[39] , \R_DATA_TEMPR84[38] , 
        \R_DATA_TEMPR84[37] , \R_DATA_TEMPR84[36] , 
        \R_DATA_TEMPR84[35] , \R_DATA_TEMPR84[34] , 
        \R_DATA_TEMPR84[33] , \R_DATA_TEMPR84[32] , 
        \R_DATA_TEMPR84[31] , \R_DATA_TEMPR84[30] , 
        \R_DATA_TEMPR84[29] , \R_DATA_TEMPR84[28] , 
        \R_DATA_TEMPR84[27] , \R_DATA_TEMPR84[26] , 
        \R_DATA_TEMPR84[25] , \R_DATA_TEMPR84[24] , 
        \R_DATA_TEMPR84[23] , \R_DATA_TEMPR84[22] , 
        \R_DATA_TEMPR84[21] , \R_DATA_TEMPR84[20] }), .B_DOUT({
        \R_DATA_TEMPR84[19] , \R_DATA_TEMPR84[18] , 
        \R_DATA_TEMPR84[17] , \R_DATA_TEMPR84[16] , 
        \R_DATA_TEMPR84[15] , \R_DATA_TEMPR84[14] , 
        \R_DATA_TEMPR84[13] , \R_DATA_TEMPR84[12] , 
        \R_DATA_TEMPR84[11] , \R_DATA_TEMPR84[10] , 
        \R_DATA_TEMPR84[9] , \R_DATA_TEMPR84[8] , \R_DATA_TEMPR84[7] , 
        \R_DATA_TEMPR84[6] , \R_DATA_TEMPR84[5] , \R_DATA_TEMPR84[4] , 
        \R_DATA_TEMPR84[3] , \R_DATA_TEMPR84[2] , \R_DATA_TEMPR84[1] , 
        \R_DATA_TEMPR84[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[84][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[21] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[21] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_236 (.A(\R_DATA_TEMPR8[23] ), .B(\R_DATA_TEMPR9[23] ), .C(
        \R_DATA_TEMPR10[23] ), .D(\R_DATA_TEMPR11[23] ), .Y(OR4_236_Y));
    OR4 OR4_1226 (.A(\R_DATA_TEMPR96[37] ), .B(\R_DATA_TEMPR97[37] ), 
        .C(\R_DATA_TEMPR98[37] ), .D(\R_DATA_TEMPR99[37] ), .Y(
        OR4_1226_Y));
    OR2 OR2_7 (.A(\R_DATA_TEMPR84[28] ), .B(\R_DATA_TEMPR85[28] ), .Y(
        OR2_7_Y));
    OR4 OR4_1399 (.A(OR4_282_Y), .B(OR2_20_Y), .C(\R_DATA_TEMPR86[0] ), 
        .D(\R_DATA_TEMPR87[0] ), .Y(OR4_1399_Y));
    OR4 OR4_73 (.A(\R_DATA_TEMPR40[29] ), .B(\R_DATA_TEMPR41[29] ), .C(
        \R_DATA_TEMPR42[29] ), .D(\R_DATA_TEMPR43[29] ), .Y(OR4_73_Y));
    OR4 OR4_1042 (.A(\R_DATA_TEMPR116[29] ), .B(\R_DATA_TEMPR117[29] ), 
        .C(\R_DATA_TEMPR118[29] ), .D(\R_DATA_TEMPR119[29] ), .Y(
        OR4_1042_Y));
    OR4 OR4_195 (.A(\R_DATA_TEMPR60[35] ), .B(\R_DATA_TEMPR61[35] ), 
        .C(\R_DATA_TEMPR62[35] ), .D(\R_DATA_TEMPR63[35] ), .Y(
        OR4_195_Y));
    OR4 OR4_1458 (.A(\R_DATA_TEMPR16[38] ), .B(\R_DATA_TEMPR17[38] ), 
        .C(\R_DATA_TEMPR18[38] ), .D(\R_DATA_TEMPR19[38] ), .Y(
        OR4_1458_Y));
    OR4 OR4_252 (.A(OR4_1585_Y), .B(OR4_407_Y), .C(OR4_1377_Y), .D(
        OR4_40_Y), .Y(OR4_252_Y));
    OR4 OR4_1090 (.A(\R_DATA_TEMPR40[4] ), .B(\R_DATA_TEMPR41[4] ), .C(
        \R_DATA_TEMPR42[4] ), .D(\R_DATA_TEMPR43[4] ), .Y(OR4_1090_Y));
    OR4 OR4_1328 (.A(\R_DATA_TEMPR56[18] ), .B(\R_DATA_TEMPR57[18] ), 
        .C(\R_DATA_TEMPR58[18] ), .D(\R_DATA_TEMPR59[18] ), .Y(
        OR4_1328_Y));
    OR4 OR4_289 (.A(\R_DATA_TEMPR60[9] ), .B(\R_DATA_TEMPR61[9] ), .C(
        \R_DATA_TEMPR62[9] ), .D(\R_DATA_TEMPR63[9] ), .Y(OR4_289_Y));
    OR4 OR4_1003 (.A(\R_DATA_TEMPR52[36] ), .B(\R_DATA_TEMPR53[36] ), 
        .C(\R_DATA_TEMPR54[36] ), .D(\R_DATA_TEMPR55[36] ), .Y(
        OR4_1003_Y));
    OR4 OR4_907 (.A(OR4_1361_Y), .B(OR4_32_Y), .C(OR4_281_Y), .D(
        OR4_89_Y), .Y(OR4_907_Y));
    OR4 OR4_497 (.A(OR4_434_Y), .B(OR4_1286_Y), .C(OR4_457_Y), .D(
        OR4_706_Y), .Y(OR4_497_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%52%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R52C0 (.A_DOUT({
        \R_DATA_TEMPR52[39] , \R_DATA_TEMPR52[38] , 
        \R_DATA_TEMPR52[37] , \R_DATA_TEMPR52[36] , 
        \R_DATA_TEMPR52[35] , \R_DATA_TEMPR52[34] , 
        \R_DATA_TEMPR52[33] , \R_DATA_TEMPR52[32] , 
        \R_DATA_TEMPR52[31] , \R_DATA_TEMPR52[30] , 
        \R_DATA_TEMPR52[29] , \R_DATA_TEMPR52[28] , 
        \R_DATA_TEMPR52[27] , \R_DATA_TEMPR52[26] , 
        \R_DATA_TEMPR52[25] , \R_DATA_TEMPR52[24] , 
        \R_DATA_TEMPR52[23] , \R_DATA_TEMPR52[22] , 
        \R_DATA_TEMPR52[21] , \R_DATA_TEMPR52[20] }), .B_DOUT({
        \R_DATA_TEMPR52[19] , \R_DATA_TEMPR52[18] , 
        \R_DATA_TEMPR52[17] , \R_DATA_TEMPR52[16] , 
        \R_DATA_TEMPR52[15] , \R_DATA_TEMPR52[14] , 
        \R_DATA_TEMPR52[13] , \R_DATA_TEMPR52[12] , 
        \R_DATA_TEMPR52[11] , \R_DATA_TEMPR52[10] , 
        \R_DATA_TEMPR52[9] , \R_DATA_TEMPR52[8] , \R_DATA_TEMPR52[7] , 
        \R_DATA_TEMPR52[6] , \R_DATA_TEMPR52[5] , \R_DATA_TEMPR52[4] , 
        \R_DATA_TEMPR52[3] , \R_DATA_TEMPR52[2] , \R_DATA_TEMPR52[1] , 
        \R_DATA_TEMPR52[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[52][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[13] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[13] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_32 (.A(\R_DATA_TEMPR84[34] ), .B(\R_DATA_TEMPR85[34] ), .Y(
        OR2_32_Y));
    OR4 OR4_634 (.A(\R_DATA_TEMPR0[10] ), .B(\R_DATA_TEMPR1[10] ), .C(
        \R_DATA_TEMPR2[10] ), .D(\R_DATA_TEMPR3[10] ), .Y(OR4_634_Y));
    OR4 OR4_1402 (.A(\R_DATA_TEMPR108[36] ), .B(\R_DATA_TEMPR109[36] ), 
        .C(\R_DATA_TEMPR110[36] ), .D(\R_DATA_TEMPR111[36] ), .Y(
        OR4_1402_Y));
    OR4 OR4_1185 (.A(OR4_590_Y), .B(OR4_416_Y), .C(OR4_1457_Y), .D(
        OR4_344_Y), .Y(OR4_1185_Y));
    OR2 OR2_1 (.A(\R_DATA_TEMPR84[4] ), .B(\R_DATA_TEMPR85[4] ), .Y(
        OR2_1_Y));
    OR4 OR4_464 (.A(\R_DATA_TEMPR108[18] ), .B(\R_DATA_TEMPR109[18] ), 
        .C(\R_DATA_TEMPR110[18] ), .D(\R_DATA_TEMPR111[18] ), .Y(
        OR4_464_Y));
    OR4 OR4_977 (.A(\R_DATA_TEMPR36[9] ), .B(\R_DATA_TEMPR37[9] ), .C(
        \R_DATA_TEMPR38[9] ), .D(\R_DATA_TEMPR39[9] ), .Y(OR4_977_Y));
    OR4 OR4_1081 (.A(\R_DATA_TEMPR88[19] ), .B(\R_DATA_TEMPR89[19] ), 
        .C(\R_DATA_TEMPR90[19] ), .D(\R_DATA_TEMPR91[19] ), .Y(
        OR4_1081_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%42%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R42C0 (.A_DOUT({
        \R_DATA_TEMPR42[39] , \R_DATA_TEMPR42[38] , 
        \R_DATA_TEMPR42[37] , \R_DATA_TEMPR42[36] , 
        \R_DATA_TEMPR42[35] , \R_DATA_TEMPR42[34] , 
        \R_DATA_TEMPR42[33] , \R_DATA_TEMPR42[32] , 
        \R_DATA_TEMPR42[31] , \R_DATA_TEMPR42[30] , 
        \R_DATA_TEMPR42[29] , \R_DATA_TEMPR42[28] , 
        \R_DATA_TEMPR42[27] , \R_DATA_TEMPR42[26] , 
        \R_DATA_TEMPR42[25] , \R_DATA_TEMPR42[24] , 
        \R_DATA_TEMPR42[23] , \R_DATA_TEMPR42[22] , 
        \R_DATA_TEMPR42[21] , \R_DATA_TEMPR42[20] }), .B_DOUT({
        \R_DATA_TEMPR42[19] , \R_DATA_TEMPR42[18] , 
        \R_DATA_TEMPR42[17] , \R_DATA_TEMPR42[16] , 
        \R_DATA_TEMPR42[15] , \R_DATA_TEMPR42[14] , 
        \R_DATA_TEMPR42[13] , \R_DATA_TEMPR42[12] , 
        \R_DATA_TEMPR42[11] , \R_DATA_TEMPR42[10] , 
        \R_DATA_TEMPR42[9] , \R_DATA_TEMPR42[8] , \R_DATA_TEMPR42[7] , 
        \R_DATA_TEMPR42[6] , \R_DATA_TEMPR42[5] , \R_DATA_TEMPR42[4] , 
        \R_DATA_TEMPR42[3] , \R_DATA_TEMPR42[2] , \R_DATA_TEMPR42[1] , 
        \R_DATA_TEMPR42[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[42][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[10] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[10] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%96%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R96C0 (.A_DOUT({
        \R_DATA_TEMPR96[39] , \R_DATA_TEMPR96[38] , 
        \R_DATA_TEMPR96[37] , \R_DATA_TEMPR96[36] , 
        \R_DATA_TEMPR96[35] , \R_DATA_TEMPR96[34] , 
        \R_DATA_TEMPR96[33] , \R_DATA_TEMPR96[32] , 
        \R_DATA_TEMPR96[31] , \R_DATA_TEMPR96[30] , 
        \R_DATA_TEMPR96[29] , \R_DATA_TEMPR96[28] , 
        \R_DATA_TEMPR96[27] , \R_DATA_TEMPR96[26] , 
        \R_DATA_TEMPR96[25] , \R_DATA_TEMPR96[24] , 
        \R_DATA_TEMPR96[23] , \R_DATA_TEMPR96[22] , 
        \R_DATA_TEMPR96[21] , \R_DATA_TEMPR96[20] }), .B_DOUT({
        \R_DATA_TEMPR96[19] , \R_DATA_TEMPR96[18] , 
        \R_DATA_TEMPR96[17] , \R_DATA_TEMPR96[16] , 
        \R_DATA_TEMPR96[15] , \R_DATA_TEMPR96[14] , 
        \R_DATA_TEMPR96[13] , \R_DATA_TEMPR96[12] , 
        \R_DATA_TEMPR96[11] , \R_DATA_TEMPR96[10] , 
        \R_DATA_TEMPR96[9] , \R_DATA_TEMPR96[8] , \R_DATA_TEMPR96[7] , 
        \R_DATA_TEMPR96[6] , \R_DATA_TEMPR96[5] , \R_DATA_TEMPR96[4] , 
        \R_DATA_TEMPR96[3] , \R_DATA_TEMPR96[2] , \R_DATA_TEMPR96[1] , 
        \R_DATA_TEMPR96[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[96][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[24] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[24] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_210 (.A(\R_DATA_TEMPR32[10] ), .B(\R_DATA_TEMPR33[10] ), 
        .C(\R_DATA_TEMPR34[10] ), .D(\R_DATA_TEMPR35[10] ), .Y(
        OR4_210_Y));
    OR4 OR4_742 (.A(\R_DATA_TEMPR16[16] ), .B(\R_DATA_TEMPR17[16] ), 
        .C(\R_DATA_TEMPR18[16] ), .D(\R_DATA_TEMPR19[16] ), .Y(
        OR4_742_Y));
    OR4 OR4_517 (.A(OR4_1426_Y), .B(OR2_14_Y), .C(\R_DATA_TEMPR86[14] )
        , .D(\R_DATA_TEMPR87[14] ), .Y(OR4_517_Y));
    OR4 OR4_350 (.A(\R_DATA_TEMPR104[9] ), .B(\R_DATA_TEMPR105[9] ), 
        .C(\R_DATA_TEMPR106[9] ), .D(\R_DATA_TEMPR107[9] ), .Y(
        OR4_350_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[1]  (.A(CFG3_8_Y), .B(CFG3_12_Y)
        , .Y(\BLKX2[1] ));
    OR4 OR4_366 (.A(\R_DATA_TEMPR112[9] ), .B(\R_DATA_TEMPR113[9] ), 
        .C(\R_DATA_TEMPR114[9] ), .D(\R_DATA_TEMPR115[9] ), .Y(
        OR4_366_Y));
    OR4 OR4_1499 (.A(OR4_448_Y), .B(OR4_986_Y), .C(OR4_1527_Y), .D(
        OR4_362_Y), .Y(OR4_1499_Y));
    OR4 OR4_295 (.A(OR4_523_Y), .B(OR4_775_Y), .C(OR4_956_Y), .D(
        OR4_1194_Y), .Y(OR4_295_Y));
    OR4 OR4_946 (.A(\R_DATA_TEMPR104[28] ), .B(\R_DATA_TEMPR105[28] ), 
        .C(\R_DATA_TEMPR106[28] ), .D(\R_DATA_TEMPR107[28] ), .Y(
        OR4_946_Y));
    OR4 OR4_1154 (.A(OR4_338_Y), .B(OR4_424_Y), .C(OR4_950_Y), .D(
        OR4_1417_Y), .Y(OR4_1154_Y));
    OR4 OR4_889 (.A(\R_DATA_TEMPR76[29] ), .B(\R_DATA_TEMPR77[29] ), 
        .C(\R_DATA_TEMPR78[29] ), .D(\R_DATA_TEMPR79[29] ), .Y(
        OR4_889_Y));
    OR4 OR4_1460 (.A(\R_DATA_TEMPR48[24] ), .B(\R_DATA_TEMPR49[24] ), 
        .C(\R_DATA_TEMPR50[24] ), .D(\R_DATA_TEMPR51[24] ), .Y(
        OR4_1460_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[17]  (.A(CFG3_15_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[17] ));
    OR4 OR4_892 (.A(\R_DATA_TEMPR96[31] ), .B(\R_DATA_TEMPR97[31] ), 
        .C(\R_DATA_TEMPR98[31] ), .D(\R_DATA_TEMPR99[31] ), .Y(
        OR4_892_Y));
    OR4 OR4_1029 (.A(OR4_622_Y), .B(OR4_923_Y), .C(OR4_382_Y), .D(
        OR4_1230_Y), .Y(OR4_1029_Y));
    OR4 OR4_645 (.A(\R_DATA_TEMPR112[39] ), .B(\R_DATA_TEMPR113[39] ), 
        .C(\R_DATA_TEMPR114[39] ), .D(\R_DATA_TEMPR115[39] ), .Y(
        OR4_645_Y));
    OR4 OR4_619 (.A(\R_DATA_TEMPR44[25] ), .B(\R_DATA_TEMPR45[25] ), 
        .C(\R_DATA_TEMPR46[25] ), .D(\R_DATA_TEMPR47[25] ), .Y(
        OR4_619_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[18]  (.A(CFG3_14_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[18] ));
    OR4 OR4_1110 (.A(\R_DATA_TEMPR36[1] ), .B(\R_DATA_TEMPR37[1] ), .C(
        \R_DATA_TEMPR38[1] ), .D(\R_DATA_TEMPR39[1] ), .Y(OR4_1110_Y));
    OR4 OR4_853 (.A(\R_DATA_TEMPR0[30] ), .B(\R_DATA_TEMPR1[30] ), .C(
        \R_DATA_TEMPR2[30] ), .D(\R_DATA_TEMPR3[30] ), .Y(OR4_853_Y));
    OR4 OR4_1083 (.A(\R_DATA_TEMPR16[34] ), .B(\R_DATA_TEMPR17[34] ), 
        .C(\R_DATA_TEMPR18[34] ), .D(\R_DATA_TEMPR19[34] ), .Y(
        OR4_1083_Y));
    OR4 OR4_1550 (.A(OR4_932_Y), .B(OR4_618_Y), .C(OR4_1034_Y), .D(
        OR4_873_Y), .Y(OR4_1550_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[13]  (.A(CFG3_22_Y), .B(
        CFG3_4_Y), .Y(\BLKX2[13] ));
    OR4 OR4_35 (.A(\R_DATA_TEMPR76[11] ), .B(\R_DATA_TEMPR77[11] ), .C(
        \R_DATA_TEMPR78[11] ), .D(\R_DATA_TEMPR79[11] ), .Y(OR4_35_Y));
    OR4 OR4_1482 (.A(\R_DATA_TEMPR120[10] ), .B(\R_DATA_TEMPR121[10] ), 
        .C(\R_DATA_TEMPR122[10] ), .D(\R_DATA_TEMPR123[10] ), .Y(
        OR4_1482_Y));
    OR4 OR4_1161 (.A(\R_DATA_TEMPR56[24] ), .B(\R_DATA_TEMPR57[24] ), 
        .C(\R_DATA_TEMPR58[24] ), .D(\R_DATA_TEMPR59[24] ), .Y(
        OR4_1161_Y));
    OR4 OR4_405 (.A(\R_DATA_TEMPR4[24] ), .B(\R_DATA_TEMPR5[24] ), .C(
        \R_DATA_TEMPR6[24] ), .D(\R_DATA_TEMPR7[24] ), .Y(OR4_405_Y));
    OR4 OR4_216 (.A(\R_DATA_TEMPR80[20] ), .B(\R_DATA_TEMPR81[20] ), 
        .C(\R_DATA_TEMPR82[20] ), .D(\R_DATA_TEMPR83[20] ), .Y(
        OR4_216_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%70%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R70C0 (.A_DOUT({
        \R_DATA_TEMPR70[39] , \R_DATA_TEMPR70[38] , 
        \R_DATA_TEMPR70[37] , \R_DATA_TEMPR70[36] , 
        \R_DATA_TEMPR70[35] , \R_DATA_TEMPR70[34] , 
        \R_DATA_TEMPR70[33] , \R_DATA_TEMPR70[32] , 
        \R_DATA_TEMPR70[31] , \R_DATA_TEMPR70[30] , 
        \R_DATA_TEMPR70[29] , \R_DATA_TEMPR70[28] , 
        \R_DATA_TEMPR70[27] , \R_DATA_TEMPR70[26] , 
        \R_DATA_TEMPR70[25] , \R_DATA_TEMPR70[24] , 
        \R_DATA_TEMPR70[23] , \R_DATA_TEMPR70[22] , 
        \R_DATA_TEMPR70[21] , \R_DATA_TEMPR70[20] }), .B_DOUT({
        \R_DATA_TEMPR70[19] , \R_DATA_TEMPR70[18] , 
        \R_DATA_TEMPR70[17] , \R_DATA_TEMPR70[16] , 
        \R_DATA_TEMPR70[15] , \R_DATA_TEMPR70[14] , 
        \R_DATA_TEMPR70[13] , \R_DATA_TEMPR70[12] , 
        \R_DATA_TEMPR70[11] , \R_DATA_TEMPR70[10] , 
        \R_DATA_TEMPR70[9] , \R_DATA_TEMPR70[8] , \R_DATA_TEMPR70[7] , 
        \R_DATA_TEMPR70[6] , \R_DATA_TEMPR70[5] , \R_DATA_TEMPR70[4] , 
        \R_DATA_TEMPR70[3] , \R_DATA_TEMPR70[2] , \R_DATA_TEMPR70[1] , 
        \R_DATA_TEMPR70[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[70][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[17] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[17] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_71 (.A(\R_DATA_TEMPR36[32] ), .B(\R_DATA_TEMPR37[32] ), .C(
        \R_DATA_TEMPR38[32] ), .D(\R_DATA_TEMPR39[32] ), .Y(OR4_71_Y));
    OR4 OR4_1258 (.A(\R_DATA_TEMPR64[2] ), .B(\R_DATA_TEMPR65[2] ), .C(
        \R_DATA_TEMPR66[2] ), .D(\R_DATA_TEMPR67[2] ), .Y(OR4_1258_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%101%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R101C0 (.A_DOUT({
        \R_DATA_TEMPR101[39] , \R_DATA_TEMPR101[38] , 
        \R_DATA_TEMPR101[37] , \R_DATA_TEMPR101[36] , 
        \R_DATA_TEMPR101[35] , \R_DATA_TEMPR101[34] , 
        \R_DATA_TEMPR101[33] , \R_DATA_TEMPR101[32] , 
        \R_DATA_TEMPR101[31] , \R_DATA_TEMPR101[30] , 
        \R_DATA_TEMPR101[29] , \R_DATA_TEMPR101[28] , 
        \R_DATA_TEMPR101[27] , \R_DATA_TEMPR101[26] , 
        \R_DATA_TEMPR101[25] , \R_DATA_TEMPR101[24] , 
        \R_DATA_TEMPR101[23] , \R_DATA_TEMPR101[22] , 
        \R_DATA_TEMPR101[21] , \R_DATA_TEMPR101[20] }), .B_DOUT({
        \R_DATA_TEMPR101[19] , \R_DATA_TEMPR101[18] , 
        \R_DATA_TEMPR101[17] , \R_DATA_TEMPR101[16] , 
        \R_DATA_TEMPR101[15] , \R_DATA_TEMPR101[14] , 
        \R_DATA_TEMPR101[13] , \R_DATA_TEMPR101[12] , 
        \R_DATA_TEMPR101[11] , \R_DATA_TEMPR101[10] , 
        \R_DATA_TEMPR101[9] , \R_DATA_TEMPR101[8] , 
        \R_DATA_TEMPR101[7] , \R_DATA_TEMPR101[6] , 
        \R_DATA_TEMPR101[5] , \R_DATA_TEMPR101[4] , 
        \R_DATA_TEMPR101[3] , \R_DATA_TEMPR101[2] , 
        \R_DATA_TEMPR101[1] , \R_DATA_TEMPR101[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[101][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[25] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[25] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_475 (.A(\R_DATA_TEMPR64[16] ), .B(\R_DATA_TEMPR65[16] ), 
        .C(\R_DATA_TEMPR66[16] ), .D(\R_DATA_TEMPR67[16] ), .Y(
        OR4_475_Y));
    OR4 OR4_1566 (.A(OR4_257_Y), .B(OR4_1318_Y), .C(OR4_1283_Y), .D(
        OR4_963_Y), .Y(OR4_1566_Y));
    OR4 OR4_125 (.A(\R_DATA_TEMPR120[11] ), .B(\R_DATA_TEMPR121[11] ), 
        .C(\R_DATA_TEMPR122[11] ), .D(\R_DATA_TEMPR123[11] ), .Y(
        OR4_125_Y));
    OR4 OR4_1543 (.A(OR4_180_Y), .B(OR4_759_Y), .C(OR4_1542_Y), .D(
        OR4_166_Y), .Y(OR4_1543_Y));
    OR4 OR4_493 (.A(\R_DATA_TEMPR60[11] ), .B(\R_DATA_TEMPR61[11] ), 
        .C(\R_DATA_TEMPR62[11] ), .D(\R_DATA_TEMPR63[11] ), .Y(
        OR4_493_Y));
    OR4 OR4_1137 (.A(\R_DATA_TEMPR72[22] ), .B(\R_DATA_TEMPR73[22] ), 
        .C(\R_DATA_TEMPR74[22] ), .D(\R_DATA_TEMPR75[22] ), .Y(
        OR4_1137_Y));
    OR4 OR4_691 (.A(OR4_165_Y), .B(OR4_1060_Y), .C(OR4_1612_Y), .D(
        OR4_995_Y), .Y(OR4_691_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%80%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R80C0 (.A_DOUT({
        \R_DATA_TEMPR80[39] , \R_DATA_TEMPR80[38] , 
        \R_DATA_TEMPR80[37] , \R_DATA_TEMPR80[36] , 
        \R_DATA_TEMPR80[35] , \R_DATA_TEMPR80[34] , 
        \R_DATA_TEMPR80[33] , \R_DATA_TEMPR80[32] , 
        \R_DATA_TEMPR80[31] , \R_DATA_TEMPR80[30] , 
        \R_DATA_TEMPR80[29] , \R_DATA_TEMPR80[28] , 
        \R_DATA_TEMPR80[27] , \R_DATA_TEMPR80[26] , 
        \R_DATA_TEMPR80[25] , \R_DATA_TEMPR80[24] , 
        \R_DATA_TEMPR80[23] , \R_DATA_TEMPR80[22] , 
        \R_DATA_TEMPR80[21] , \R_DATA_TEMPR80[20] }), .B_DOUT({
        \R_DATA_TEMPR80[19] , \R_DATA_TEMPR80[18] , 
        \R_DATA_TEMPR80[17] , \R_DATA_TEMPR80[16] , 
        \R_DATA_TEMPR80[15] , \R_DATA_TEMPR80[14] , 
        \R_DATA_TEMPR80[13] , \R_DATA_TEMPR80[12] , 
        \R_DATA_TEMPR80[11] , \R_DATA_TEMPR80[10] , 
        \R_DATA_TEMPR80[9] , \R_DATA_TEMPR80[8] , \R_DATA_TEMPR80[7] , 
        \R_DATA_TEMPR80[6] , \R_DATA_TEMPR80[5] , \R_DATA_TEMPR80[4] , 
        \R_DATA_TEMPR80[3] , \R_DATA_TEMPR80[2] , \R_DATA_TEMPR80[1] , 
        \R_DATA_TEMPR80[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[80][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[20] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[20] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_614 (.A(\R_DATA_TEMPR56[33] ), .B(\R_DATA_TEMPR57[33] ), 
        .C(\R_DATA_TEMPR58[33] ), .D(\R_DATA_TEMPR59[33] ), .Y(
        OR4_614_Y));
    OR4 OR4_427 (.A(OR4_1584_Y), .B(OR4_973_Y), .C(OR4_1220_Y), .D(
        OR4_160_Y), .Y(OR4_427_Y));
    OR4 OR4_1008 (.A(\R_DATA_TEMPR120[30] ), .B(\R_DATA_TEMPR121[30] ), 
        .C(\R_DATA_TEMPR122[30] ), .D(\R_DATA_TEMPR123[30] ), .Y(
        OR4_1008_Y));
    OR4 OR4_787 (.A(OR4_301_Y), .B(OR4_640_Y), .C(OR4_610_Y), .D(
        OR4_1408_Y), .Y(OR4_787_Y));
    OR4 OR4_298 (.A(\R_DATA_TEMPR52[29] ), .B(\R_DATA_TEMPR53[29] ), 
        .C(\R_DATA_TEMPR54[29] ), .D(\R_DATA_TEMPR55[29] ), .Y(
        OR4_298_Y));
    OR4 \OR4_R_DATA[27]  (.A(OR4_215_Y), .B(OR4_988_Y), .C(OR4_1421_Y), 
        .D(OR4_1563_Y), .Y(R_DATA[27]));
    OR4 OR4_784 (.A(\R_DATA_TEMPR20[39] ), .B(\R_DATA_TEMPR21[39] ), 
        .C(\R_DATA_TEMPR22[39] ), .D(\R_DATA_TEMPR23[39] ), .Y(
        OR4_784_Y));
    OR4 OR4_1310 (.A(\R_DATA_TEMPR64[23] ), .B(\R_DATA_TEMPR65[23] ), 
        .C(\R_DATA_TEMPR66[23] ), .D(\R_DATA_TEMPR67[23] ), .Y(
        OR4_1310_Y));
    OR4 OR4_28 (.A(OR4_119_Y), .B(OR4_1452_Y), .C(OR4_233_Y), .D(
        OR4_58_Y), .Y(OR4_28_Y));
    OR4 OR4_1277 (.A(\R_DATA_TEMPR124[29] ), .B(\R_DATA_TEMPR125[29] ), 
        .C(\R_DATA_TEMPR126[29] ), .D(\R_DATA_TEMPR127[29] ), .Y(
        OR4_1277_Y));
    OR4 OR4_640 (.A(\R_DATA_TEMPR36[19] ), .B(\R_DATA_TEMPR37[19] ), 
        .C(\R_DATA_TEMPR38[19] ), .D(\R_DATA_TEMPR39[19] ), .Y(
        OR4_640_Y));
    OR4 OR4_881 (.A(\R_DATA_TEMPR8[9] ), .B(\R_DATA_TEMPR9[9] ), .C(
        \R_DATA_TEMPR10[9] ), .D(\R_DATA_TEMPR11[9] ), .Y(OR4_881_Y));
    OR4 OR4_1502 (.A(OR4_472_Y), .B(OR4_915_Y), .C(OR4_259_Y), .D(
        OR4_567_Y), .Y(OR4_1502_Y));
    OR4 OR4_1490 (.A(\R_DATA_TEMPR32[39] ), .B(\R_DATA_TEMPR33[39] ), 
        .C(\R_DATA_TEMPR34[39] ), .D(\R_DATA_TEMPR35[39] ), .Y(
        OR4_1490_Y));
    OR4 OR4_1467 (.A(\R_DATA_TEMPR8[35] ), .B(\R_DATA_TEMPR9[35] ), .C(
        \R_DATA_TEMPR10[35] ), .D(\R_DATA_TEMPR11[35] ), .Y(OR4_1467_Y)
        );
    OR4 OR4_164 (.A(\R_DATA_TEMPR40[24] ), .B(\R_DATA_TEMPR41[24] ), 
        .C(\R_DATA_TEMPR42[24] ), .D(\R_DATA_TEMPR43[24] ), .Y(
        OR4_164_Y));
    OR4 OR4_404 (.A(\R_DATA_TEMPR112[5] ), .B(\R_DATA_TEMPR113[5] ), 
        .C(\R_DATA_TEMPR114[5] ), .D(\R_DATA_TEMPR115[5] ), .Y(
        OR4_404_Y));
    OR4 OR4_225 (.A(\R_DATA_TEMPR20[23] ), .B(\R_DATA_TEMPR21[23] ), 
        .C(\R_DATA_TEMPR22[23] ), .D(\R_DATA_TEMPR23[23] ), .Y(
        OR4_225_Y));
    OR4 OR4_555 (.A(\R_DATA_TEMPR20[16] ), .B(\R_DATA_TEMPR21[16] ), 
        .C(\R_DATA_TEMPR22[16] ), .D(\R_DATA_TEMPR23[16] ), .Y(
        OR4_555_Y));
    OR4 OR4_347 (.A(\R_DATA_TEMPR80[19] ), .B(\R_DATA_TEMPR81[19] ), 
        .C(\R_DATA_TEMPR82[19] ), .D(\R_DATA_TEMPR83[19] ), .Y(
        OR4_347_Y));
    OR4 OR4_140 (.A(\R_DATA_TEMPR48[32] ), .B(\R_DATA_TEMPR49[32] ), 
        .C(\R_DATA_TEMPR50[32] ), .D(\R_DATA_TEMPR51[32] ), .Y(
        OR4_140_Y));
    OR4 OR4_822 (.A(\R_DATA_TEMPR124[28] ), .B(\R_DATA_TEMPR125[28] ), 
        .C(\R_DATA_TEMPR126[28] ), .D(\R_DATA_TEMPR127[28] ), .Y(
        OR4_822_Y));
    OR4 OR4_1476 (.A(\R_DATA_TEMPR104[0] ), .B(\R_DATA_TEMPR105[0] ), 
        .C(\R_DATA_TEMPR106[0] ), .D(\R_DATA_TEMPR107[0] ), .Y(
        OR4_1476_Y));
    OR4 OR4_1374 (.A(\R_DATA_TEMPR40[38] ), .B(\R_DATA_TEMPR41[38] ), 
        .C(\R_DATA_TEMPR42[38] ), .D(\R_DATA_TEMPR43[38] ), .Y(
        OR4_1374_Y));
    OR4 OR4_1065 (.A(\R_DATA_TEMPR104[17] ), .B(\R_DATA_TEMPR105[17] ), 
        .C(\R_DATA_TEMPR106[17] ), .D(\R_DATA_TEMPR107[17] ), .Y(
        OR4_1065_Y));
    OR4 OR4_474 (.A(\R_DATA_TEMPR4[36] ), .B(\R_DATA_TEMPR5[36] ), .C(
        \R_DATA_TEMPR6[36] ), .D(\R_DATA_TEMPR7[36] ), .Y(OR4_474_Y));
    OR4 OR4_1191 (.A(\R_DATA_TEMPR44[24] ), .B(\R_DATA_TEMPR45[24] ), 
        .C(\R_DATA_TEMPR46[24] ), .D(\R_DATA_TEMPR47[24] ), .Y(
        OR4_1191_Y));
    OR4 OR4_306 (.A(OR4_786_Y), .B(OR4_474_Y), .C(OR4_902_Y), .D(
        OR4_720_Y), .Y(OR4_306_Y));
    OR4 OR4_1088 (.A(OR4_1458_Y), .B(OR4_346_Y), .C(OR4_1480_Y), .D(
        OR4_965_Y), .Y(OR4_1088_Y));
    OR4 OR4_963 (.A(\R_DATA_TEMPR44[33] ), .B(\R_DATA_TEMPR45[33] ), 
        .C(\R_DATA_TEMPR46[33] ), .D(\R_DATA_TEMPR47[33] ), .Y(
        OR4_963_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%124%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R124C0 (.A_DOUT({
        \R_DATA_TEMPR124[39] , \R_DATA_TEMPR124[38] , 
        \R_DATA_TEMPR124[37] , \R_DATA_TEMPR124[36] , 
        \R_DATA_TEMPR124[35] , \R_DATA_TEMPR124[34] , 
        \R_DATA_TEMPR124[33] , \R_DATA_TEMPR124[32] , 
        \R_DATA_TEMPR124[31] , \R_DATA_TEMPR124[30] , 
        \R_DATA_TEMPR124[29] , \R_DATA_TEMPR124[28] , 
        \R_DATA_TEMPR124[27] , \R_DATA_TEMPR124[26] , 
        \R_DATA_TEMPR124[25] , \R_DATA_TEMPR124[24] , 
        \R_DATA_TEMPR124[23] , \R_DATA_TEMPR124[22] , 
        \R_DATA_TEMPR124[21] , \R_DATA_TEMPR124[20] }), .B_DOUT({
        \R_DATA_TEMPR124[19] , \R_DATA_TEMPR124[18] , 
        \R_DATA_TEMPR124[17] , \R_DATA_TEMPR124[16] , 
        \R_DATA_TEMPR124[15] , \R_DATA_TEMPR124[14] , 
        \R_DATA_TEMPR124[13] , \R_DATA_TEMPR124[12] , 
        \R_DATA_TEMPR124[11] , \R_DATA_TEMPR124[10] , 
        \R_DATA_TEMPR124[9] , \R_DATA_TEMPR124[8] , 
        \R_DATA_TEMPR124[7] , \R_DATA_TEMPR124[6] , 
        \R_DATA_TEMPR124[5] , \R_DATA_TEMPR124[4] , 
        \R_DATA_TEMPR124[3] , \R_DATA_TEMPR124[2] , 
        \R_DATA_TEMPR124[1] , \R_DATA_TEMPR124[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[124][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[31] , \BLKY1[0] , \BLKY0[0] }), 
        .A_CLK(CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], 
        W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], 
        W_DATA[31], W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], 
        W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], 
        W_DATA[21], W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], 
        WBYTE_EN[2]}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], 
        W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], 
        W_ADDR[0], GND, GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[31] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA[19], 
        W_DATA[18], W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], 
        W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], W_DATA[9], 
        W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], 
        W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_748 (.A(\R_DATA_TEMPR96[3] ), .B(\R_DATA_TEMPR97[3] ), .C(
        \R_DATA_TEMPR98[3] ), .D(\R_DATA_TEMPR99[3] ), .Y(OR4_748_Y));
    OR4 OR4_653 (.A(OR4_636_Y), .B(OR4_128_Y), .C(OR4_193_Y), .D(
        OR4_1254_Y), .Y(OR4_653_Y));
    OR4 OR4_1155 (.A(OR4_510_Y), .B(OR4_1076_Y), .C(OR4_1619_Y), .D(
        OR4_437_Y), .Y(OR4_1155_Y));
    OR4 OR4_1596 (.A(\R_DATA_TEMPR40[30] ), .B(\R_DATA_TEMPR41[30] ), 
        .C(\R_DATA_TEMPR42[30] ), .D(\R_DATA_TEMPR43[30] ), .Y(
        OR4_1596_Y));
    OR4 OR4_376 (.A(\R_DATA_TEMPR92[34] ), .B(\R_DATA_TEMPR93[34] ), 
        .C(\R_DATA_TEMPR94[34] ), .D(\R_DATA_TEMPR95[34] ), .Y(
        OR4_376_Y));
    OR4 OR4_866 (.A(OR4_1472_Y), .B(OR4_86_Y), .C(OR4_274_Y), .D(
        OR4_1567_Y), .Y(OR4_866_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[18]  (.A(CFG3_0_Y), .B(CFG3_9_Y)
        , .Y(\BLKY2[18] ));
    OR4 OR4_1051 (.A(\R_DATA_TEMPR100[3] ), .B(\R_DATA_TEMPR101[3] ), 
        .C(\R_DATA_TEMPR102[3] ), .D(\R_DATA_TEMPR103[3] ), .Y(
        OR4_1051_Y));
    OR4 OR4_761 (.A(\R_DATA_TEMPR44[36] ), .B(\R_DATA_TEMPR45[36] ), 
        .C(\R_DATA_TEMPR46[36] ), .D(\R_DATA_TEMPR47[36] ), .Y(
        OR4_761_Y));
    OR4 OR4_1127 (.A(\R_DATA_TEMPR28[17] ), .B(\R_DATA_TEMPR29[17] ), 
        .C(\R_DATA_TEMPR30[17] ), .D(\R_DATA_TEMPR31[17] ), .Y(
        OR4_1127_Y));
    OR4 OR4_1582 (.A(OR4_1398_Y), .B(OR4_64_Y), .C(OR4_1133_Y), .D(
        OR4_371_Y), .Y(OR4_1582_Y));
    OR4 OR4_1215 (.A(\R_DATA_TEMPR68[31] ), .B(\R_DATA_TEMPR69[31] ), 
        .C(\R_DATA_TEMPR70[31] ), .D(\R_DATA_TEMPR71[31] ), .Y(
        OR4_1215_Y));
    OR4 OR4_423 (.A(\R_DATA_TEMPR48[6] ), .B(\R_DATA_TEMPR49[6] ), .C(
        \R_DATA_TEMPR50[6] ), .D(\R_DATA_TEMPR51[6] ), .Y(OR4_423_Y));
    OR4 OR4_621 (.A(\R_DATA_TEMPR104[39] ), .B(\R_DATA_TEMPR105[39] ), 
        .C(\R_DATA_TEMPR106[39] ), .D(\R_DATA_TEMPR107[39] ), .Y(
        OR4_621_Y));
    OR4 OR4_84 (.A(OR4_1587_Y), .B(OR4_1235_Y), .C(OR4_1603_Y), .D(
        OR4_702_Y), .Y(OR4_84_Y));
    OR4 OR4_1511 (.A(\R_DATA_TEMPR96[10] ), .B(\R_DATA_TEMPR97[10] ), 
        .C(\R_DATA_TEMPR98[10] ), .D(\R_DATA_TEMPR99[10] ), .Y(
        OR4_1511_Y));
    OR4 OR4_1230 (.A(\R_DATA_TEMPR108[5] ), .B(\R_DATA_TEMPR109[5] ), 
        .C(\R_DATA_TEMPR110[5] ), .D(\R_DATA_TEMPR111[5] ), .Y(
        OR4_1230_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[13]  (.A(CFG3_11_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[13] ));
    OR4 OR4_847 (.A(OR4_665_Y), .B(OR4_430_Y), .C(OR4_957_Y), .D(
        OR4_1423_Y), .Y(OR4_847_Y));
    OR4 OR4_148 (.A(\R_DATA_TEMPR72[27] ), .B(\R_DATA_TEMPR73[27] ), 
        .C(\R_DATA_TEMPR74[27] ), .D(\R_DATA_TEMPR75[27] ), .Y(
        OR4_148_Y));
    OR4 OR4_944 (.A(\R_DATA_TEMPR80[32] ), .B(\R_DATA_TEMPR81[32] ), 
        .C(\R_DATA_TEMPR82[32] ), .D(\R_DATA_TEMPR83[32] ), .Y(
        OR4_944_Y));
    OR4 OR4_228 (.A(\R_DATA_TEMPR16[17] ), .B(\R_DATA_TEMPR17[17] ), 
        .C(\R_DATA_TEMPR18[17] ), .D(\R_DATA_TEMPR19[17] ), .Y(
        OR4_228_Y));
    OR4 OR4_838 (.A(\R_DATA_TEMPR40[20] ), .B(\R_DATA_TEMPR41[20] ), 
        .C(\R_DATA_TEMPR42[20] ), .D(\R_DATA_TEMPR43[20] ), .Y(
        OR4_838_Y));
    OR4 OR4_1379 (.A(\R_DATA_TEMPR64[15] ), .B(\R_DATA_TEMPR65[15] ), 
        .C(\R_DATA_TEMPR66[15] ), .D(\R_DATA_TEMPR67[15] ), .Y(
        OR4_1379_Y));
    OR4 OR4_987 (.A(\R_DATA_TEMPR52[13] ), .B(\R_DATA_TEMPR53[13] ), 
        .C(\R_DATA_TEMPR54[13] ), .D(\R_DATA_TEMPR55[13] ), .Y(
        OR4_987_Y));
    OR4 OR4_959 (.A(\R_DATA_TEMPR44[27] ), .B(\R_DATA_TEMPR45[27] ), 
        .C(\R_DATA_TEMPR46[27] ), .D(\R_DATA_TEMPR47[27] ), .Y(
        OR4_959_Y));
    OR4 OR4_950 (.A(\R_DATA_TEMPR88[6] ), .B(\R_DATA_TEMPR89[6] ), .C(
        \R_DATA_TEMPR90[6] ), .D(\R_DATA_TEMPR91[6] ), .Y(OR4_950_Y));
    OR4 OR4_566 (.A(\R_DATA_TEMPR12[10] ), .B(\R_DATA_TEMPR13[10] ), 
        .C(\R_DATA_TEMPR14[10] ), .D(\R_DATA_TEMPR15[10] ), .Y(
        OR4_566_Y));
    OR4 OR4_591 (.A(\R_DATA_TEMPR100[27] ), .B(\R_DATA_TEMPR101[27] ), 
        .C(\R_DATA_TEMPR102[27] ), .D(\R_DATA_TEMPR103[27] ), .Y(
        OR4_591_Y));
    OR4 OR4_1497 (.A(\R_DATA_TEMPR20[9] ), .B(\R_DATA_TEMPR21[9] ), .C(
        \R_DATA_TEMPR22[9] ), .D(\R_DATA_TEMPR23[9] ), .Y(OR4_1497_Y));
    OR4 OR4_1053 (.A(OR4_273_Y), .B(OR4_1043_Y), .C(OR4_1513_Y), .D(
        OR4_190_Y), .Y(OR4_1053_Y));
    CFG3 #( .INIT(8'h20) )  CFG3_4 (.A(W_EN), .B(W_ADDR[15]), .C(
        W_ADDR[14]), .Y(CFG3_4_Y));
    OR4 OR4_1537 (.A(OR4_1123_Y), .B(OR4_287_Y), .C(OR4_744_Y), .D(
        OR4_1049_Y), .Y(OR4_1537_Y));
    OR4 OR4_1070 (.A(\R_DATA_TEMPR48[3] ), .B(\R_DATA_TEMPR49[3] ), .C(
        \R_DATA_TEMPR50[3] ), .D(\R_DATA_TEMPR51[3] ), .Y(OR4_1070_Y));
    OR4 OR4_1007 (.A(\R_DATA_TEMPR80[13] ), .B(\R_DATA_TEMPR81[13] ), 
        .C(\R_DATA_TEMPR82[13] ), .D(\R_DATA_TEMPR83[13] ), .Y(
        OR4_1007_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%12%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C0 (.A_DOUT({
        \R_DATA_TEMPR12[39] , \R_DATA_TEMPR12[38] , 
        \R_DATA_TEMPR12[37] , \R_DATA_TEMPR12[36] , 
        \R_DATA_TEMPR12[35] , \R_DATA_TEMPR12[34] , 
        \R_DATA_TEMPR12[33] , \R_DATA_TEMPR12[32] , 
        \R_DATA_TEMPR12[31] , \R_DATA_TEMPR12[30] , 
        \R_DATA_TEMPR12[29] , \R_DATA_TEMPR12[28] , 
        \R_DATA_TEMPR12[27] , \R_DATA_TEMPR12[26] , 
        \R_DATA_TEMPR12[25] , \R_DATA_TEMPR12[24] , 
        \R_DATA_TEMPR12[23] , \R_DATA_TEMPR12[22] , 
        \R_DATA_TEMPR12[21] , \R_DATA_TEMPR12[20] }), .B_DOUT({
        \R_DATA_TEMPR12[19] , \R_DATA_TEMPR12[18] , 
        \R_DATA_TEMPR12[17] , \R_DATA_TEMPR12[16] , 
        \R_DATA_TEMPR12[15] , \R_DATA_TEMPR12[14] , 
        \R_DATA_TEMPR12[13] , \R_DATA_TEMPR12[12] , 
        \R_DATA_TEMPR12[11] , \R_DATA_TEMPR12[10] , 
        \R_DATA_TEMPR12[9] , \R_DATA_TEMPR12[8] , \R_DATA_TEMPR12[7] , 
        \R_DATA_TEMPR12[6] , \R_DATA_TEMPR12[5] , \R_DATA_TEMPR12[4] , 
        \R_DATA_TEMPR12[3] , \R_DATA_TEMPR12[2] , \R_DATA_TEMPR12[1] , 
        \R_DATA_TEMPR12[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[9]  (.A(CFG3_8_Y), .B(CFG3_4_Y), 
        .Y(\BLKX2[9] ));
    OR4 OR4_1452 (.A(\R_DATA_TEMPR4[34] ), .B(\R_DATA_TEMPR5[34] ), .C(
        \R_DATA_TEMPR6[34] ), .D(\R_DATA_TEMPR7[34] ), .Y(OR4_1452_Y));
    OR4 OR4_1332 (.A(\R_DATA_TEMPR88[16] ), .B(\R_DATA_TEMPR89[16] ), 
        .C(\R_DATA_TEMPR90[16] ), .D(\R_DATA_TEMPR91[16] ), .Y(
        OR4_1332_Y));
    OR4 OR4_153 (.A(\R_DATA_TEMPR100[24] ), .B(\R_DATA_TEMPR101[24] ), 
        .C(\R_DATA_TEMPR102[24] ), .D(\R_DATA_TEMPR103[24] ), .Y(
        OR4_153_Y));
    OR4 OR4_1232 (.A(\R_DATA_TEMPR120[34] ), .B(\R_DATA_TEMPR121[34] ), 
        .C(\R_DATA_TEMPR122[34] ), .D(\R_DATA_TEMPR123[34] ), .Y(
        OR4_1232_Y));
    OR4 OR4_1095 (.A(\R_DATA_TEMPR28[23] ), .B(\R_DATA_TEMPR29[23] ), 
        .C(\R_DATA_TEMPR30[23] ), .D(\R_DATA_TEMPR31[23] ), .Y(
        OR4_1095_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%3%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C0 (.A_DOUT({
        \R_DATA_TEMPR3[39] , \R_DATA_TEMPR3[38] , \R_DATA_TEMPR3[37] , 
        \R_DATA_TEMPR3[36] , \R_DATA_TEMPR3[35] , \R_DATA_TEMPR3[34] , 
        \R_DATA_TEMPR3[33] , \R_DATA_TEMPR3[32] , \R_DATA_TEMPR3[31] , 
        \R_DATA_TEMPR3[30] , \R_DATA_TEMPR3[29] , \R_DATA_TEMPR3[28] , 
        \R_DATA_TEMPR3[27] , \R_DATA_TEMPR3[26] , \R_DATA_TEMPR3[25] , 
        \R_DATA_TEMPR3[24] , \R_DATA_TEMPR3[23] , \R_DATA_TEMPR3[22] , 
        \R_DATA_TEMPR3[21] , \R_DATA_TEMPR3[20] }), .B_DOUT({
        \R_DATA_TEMPR3[19] , \R_DATA_TEMPR3[18] , \R_DATA_TEMPR3[17] , 
        \R_DATA_TEMPR3[16] , \R_DATA_TEMPR3[15] , \R_DATA_TEMPR3[14] , 
        \R_DATA_TEMPR3[13] , \R_DATA_TEMPR3[12] , \R_DATA_TEMPR3[11] , 
        \R_DATA_TEMPR3[10] , \R_DATA_TEMPR3[9] , \R_DATA_TEMPR3[8] , 
        \R_DATA_TEMPR3[7] , \R_DATA_TEMPR3[6] , \R_DATA_TEMPR3[5] , 
        \R_DATA_TEMPR3[4] , \R_DATA_TEMPR3[3] , \R_DATA_TEMPR3[2] , 
        \R_DATA_TEMPR3[1] , \R_DATA_TEMPR3[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[3][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_9 (.A(\R_DATA_TEMPR44[16] ), .B(\R_DATA_TEMPR45[16] ), .C(
        \R_DATA_TEMPR46[16] ), .D(\R_DATA_TEMPR47[16] ), .Y(OR4_9_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%123%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R123C0 (.A_DOUT({
        \R_DATA_TEMPR123[39] , \R_DATA_TEMPR123[38] , 
        \R_DATA_TEMPR123[37] , \R_DATA_TEMPR123[36] , 
        \R_DATA_TEMPR123[35] , \R_DATA_TEMPR123[34] , 
        \R_DATA_TEMPR123[33] , \R_DATA_TEMPR123[32] , 
        \R_DATA_TEMPR123[31] , \R_DATA_TEMPR123[30] , 
        \R_DATA_TEMPR123[29] , \R_DATA_TEMPR123[28] , 
        \R_DATA_TEMPR123[27] , \R_DATA_TEMPR123[26] , 
        \R_DATA_TEMPR123[25] , \R_DATA_TEMPR123[24] , 
        \R_DATA_TEMPR123[23] , \R_DATA_TEMPR123[22] , 
        \R_DATA_TEMPR123[21] , \R_DATA_TEMPR123[20] }), .B_DOUT({
        \R_DATA_TEMPR123[19] , \R_DATA_TEMPR123[18] , 
        \R_DATA_TEMPR123[17] , \R_DATA_TEMPR123[16] , 
        \R_DATA_TEMPR123[15] , \R_DATA_TEMPR123[14] , 
        \R_DATA_TEMPR123[13] , \R_DATA_TEMPR123[12] , 
        \R_DATA_TEMPR123[11] , \R_DATA_TEMPR123[10] , 
        \R_DATA_TEMPR123[9] , \R_DATA_TEMPR123[8] , 
        \R_DATA_TEMPR123[7] , \R_DATA_TEMPR123[6] , 
        \R_DATA_TEMPR123[5] , \R_DATA_TEMPR123[4] , 
        \R_DATA_TEMPR123[3] , \R_DATA_TEMPR123[2] , 
        \R_DATA_TEMPR123[1] , \R_DATA_TEMPR123[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[123][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[30] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[30] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1443 (.A(\R_DATA_TEMPR68[5] ), .B(\R_DATA_TEMPR69[5] ), .C(
        \R_DATA_TEMPR70[5] ), .D(\R_DATA_TEMPR71[5] ), .Y(OR4_1443_Y));
    OR4 OR4_231 (.A(\R_DATA_TEMPR16[12] ), .B(\R_DATA_TEMPR17[12] ), 
        .C(\R_DATA_TEMPR18[12] ), .D(\R_DATA_TEMPR19[12] ), .Y(
        OR4_231_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%78%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R78C0 (.A_DOUT({
        \R_DATA_TEMPR78[39] , \R_DATA_TEMPR78[38] , 
        \R_DATA_TEMPR78[37] , \R_DATA_TEMPR78[36] , 
        \R_DATA_TEMPR78[35] , \R_DATA_TEMPR78[34] , 
        \R_DATA_TEMPR78[33] , \R_DATA_TEMPR78[32] , 
        \R_DATA_TEMPR78[31] , \R_DATA_TEMPR78[30] , 
        \R_DATA_TEMPR78[29] , \R_DATA_TEMPR78[28] , 
        \R_DATA_TEMPR78[27] , \R_DATA_TEMPR78[26] , 
        \R_DATA_TEMPR78[25] , \R_DATA_TEMPR78[24] , 
        \R_DATA_TEMPR78[23] , \R_DATA_TEMPR78[22] , 
        \R_DATA_TEMPR78[21] , \R_DATA_TEMPR78[20] }), .B_DOUT({
        \R_DATA_TEMPR78[19] , \R_DATA_TEMPR78[18] , 
        \R_DATA_TEMPR78[17] , \R_DATA_TEMPR78[16] , 
        \R_DATA_TEMPR78[15] , \R_DATA_TEMPR78[14] , 
        \R_DATA_TEMPR78[13] , \R_DATA_TEMPR78[12] , 
        \R_DATA_TEMPR78[11] , \R_DATA_TEMPR78[10] , 
        \R_DATA_TEMPR78[9] , \R_DATA_TEMPR78[8] , \R_DATA_TEMPR78[7] , 
        \R_DATA_TEMPR78[6] , \R_DATA_TEMPR78[5] , \R_DATA_TEMPR78[4] , 
        \R_DATA_TEMPR78[3] , \R_DATA_TEMPR78[2] , \R_DATA_TEMPR78[1] , 
        \R_DATA_TEMPR78[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[78][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[19] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[19] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1434 (.A(OR4_275_Y), .B(OR4_1114_Y), .C(OR4_27_Y), .D(
        OR4_1052_Y), .Y(OR4_1434_Y));
    OR4 OR4_104 (.A(\R_DATA_TEMPR68[25] ), .B(\R_DATA_TEMPR69[25] ), 
        .C(\R_DATA_TEMPR70[25] ), .D(\R_DATA_TEMPR71[25] ), .Y(
        OR4_104_Y));
    OR4 OR4_1479 (.A(\R_DATA_TEMPR40[12] ), .B(\R_DATA_TEMPR41[12] ), 
        .C(\R_DATA_TEMPR42[12] ), .D(\R_DATA_TEMPR43[12] ), .Y(
        OR4_1479_Y));
    OR4 OR4_292 (.A(\R_DATA_TEMPR92[2] ), .B(\R_DATA_TEMPR93[2] ), .C(
        \R_DATA_TEMPR94[2] ), .D(\R_DATA_TEMPR95[2] ), .Y(OR4_292_Y));
    CFG3 #( .INIT(8'h40) )  CFG3_5 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_5_Y));
    OR4 OR4_1160 (.A(\R_DATA_TEMPR96[13] ), .B(\R_DATA_TEMPR97[13] ), 
        .C(\R_DATA_TEMPR98[13] ), .D(\R_DATA_TEMPR99[13] ), .Y(
        OR4_1160_Y));
    OR4 OR4_1234 (.A(\R_DATA_TEMPR28[3] ), .B(\R_DATA_TEMPR29[3] ), .C(
        \R_DATA_TEMPR30[3] ), .D(\R_DATA_TEMPR31[3] ), .Y(OR4_1234_Y));
    OR4 OR4_174 (.A(\R_DATA_TEMPR80[2] ), .B(\R_DATA_TEMPR81[2] ), .C(
        \R_DATA_TEMPR82[2] ), .D(\R_DATA_TEMPR83[2] ), .Y(OR4_174_Y));
    OR2 OR2_34 (.A(\R_DATA_TEMPR84[17] ), .B(\R_DATA_TEMPR85[17] ), .Y(
        OR2_34_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%88%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R88C0 (.A_DOUT({
        \R_DATA_TEMPR88[39] , \R_DATA_TEMPR88[38] , 
        \R_DATA_TEMPR88[37] , \R_DATA_TEMPR88[36] , 
        \R_DATA_TEMPR88[35] , \R_DATA_TEMPR88[34] , 
        \R_DATA_TEMPR88[33] , \R_DATA_TEMPR88[32] , 
        \R_DATA_TEMPR88[31] , \R_DATA_TEMPR88[30] , 
        \R_DATA_TEMPR88[29] , \R_DATA_TEMPR88[28] , 
        \R_DATA_TEMPR88[27] , \R_DATA_TEMPR88[26] , 
        \R_DATA_TEMPR88[25] , \R_DATA_TEMPR88[24] , 
        \R_DATA_TEMPR88[23] , \R_DATA_TEMPR88[22] , 
        \R_DATA_TEMPR88[21] , \R_DATA_TEMPR88[20] }), .B_DOUT({
        \R_DATA_TEMPR88[19] , \R_DATA_TEMPR88[18] , 
        \R_DATA_TEMPR88[17] , \R_DATA_TEMPR88[16] , 
        \R_DATA_TEMPR88[15] , \R_DATA_TEMPR88[14] , 
        \R_DATA_TEMPR88[13] , \R_DATA_TEMPR88[12] , 
        \R_DATA_TEMPR88[11] , \R_DATA_TEMPR88[10] , 
        \R_DATA_TEMPR88[9] , \R_DATA_TEMPR88[8] , \R_DATA_TEMPR88[7] , 
        \R_DATA_TEMPR88[6] , \R_DATA_TEMPR88[5] , \R_DATA_TEMPR88[4] , 
        \R_DATA_TEMPR88[3] , \R_DATA_TEMPR88[2] , \R_DATA_TEMPR88[1] , 
        \R_DATA_TEMPR88[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[88][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[22] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[22] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_485 (.A(\R_DATA_TEMPR88[30] ), .B(\R_DATA_TEMPR89[30] ), 
        .C(\R_DATA_TEMPR90[30] ), .D(\R_DATA_TEMPR91[30] ), .Y(
        OR4_485_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[29]  (.A(CFG3_22_Y), .B(
        CFG3_7_Y), .Y(\BLKX2[29] ));
    OR4 OR4_1337 (.A(\R_DATA_TEMPR56[26] ), .B(\R_DATA_TEMPR57[26] ), 
        .C(\R_DATA_TEMPR58[26] ), .D(\R_DATA_TEMPR59[26] ), .Y(
        OR4_1337_Y));
    OR4 OR4_1087 (.A(\R_DATA_TEMPR0[9] ), .B(\R_DATA_TEMPR1[9] ), .C(
        \R_DATA_TEMPR2[9] ), .D(\R_DATA_TEMPR3[9] ), .Y(OR4_1087_Y));
    OR4 OR4_903 (.A(\R_DATA_TEMPR76[1] ), .B(\R_DATA_TEMPR77[1] ), .C(
        \R_DATA_TEMPR78[1] ), .D(\R_DATA_TEMPR79[1] ), .Y(OR4_903_Y));
    OR4 OR4_568 (.A(OR4_494_Y), .B(OR4_1268_Y), .C(OR4_103_Y), .D(
        OR4_415_Y), .Y(OR4_568_Y));
    OR4 OR4_1608 (.A(\R_DATA_TEMPR16[7] ), .B(\R_DATA_TEMPR17[7] ), .C(
        \R_DATA_TEMPR18[7] ), .D(\R_DATA_TEMPR19[7] ), .Y(OR4_1608_Y));
    OR4 OR4_1220 (.A(\R_DATA_TEMPR8[21] ), .B(\R_DATA_TEMPR9[21] ), .C(
        \R_DATA_TEMPR10[21] ), .D(\R_DATA_TEMPR11[21] ), .Y(OR4_1220_Y)
        );
    OR4 OR4_532 (.A(\R_DATA_TEMPR12[7] ), .B(\R_DATA_TEMPR13[7] ), .C(
        \R_DATA_TEMPR14[7] ), .D(\R_DATA_TEMPR15[7] ), .Y(OR4_532_Y));
    OR4 OR4_56 (.A(\R_DATA_TEMPR52[15] ), .B(\R_DATA_TEMPR53[15] ), .C(
        \R_DATA_TEMPR54[15] ), .D(\R_DATA_TEMPR55[15] ), .Y(OR4_56_Y));
    OR4 OR4_1616 (.A(\R_DATA_TEMPR52[32] ), .B(\R_DATA_TEMPR53[32] ), 
        .C(\R_DATA_TEMPR54[32] ), .D(\R_DATA_TEMPR55[32] ), .Y(
        OR4_1616_Y));
    OR4 OR4_390 (.A(OR4_1030_Y), .B(OR4_1588_Y), .C(OR4_656_Y), .D(
        OR4_1329_Y), .Y(OR4_390_Y));
    OR4 OR4_818 (.A(OR4_252_Y), .B(OR4_356_Y), .C(OR4_877_Y), .D(
        OR4_343_Y), .Y(OR4_818_Y));
    OR4 OR4_973 (.A(\R_DATA_TEMPR4[21] ), .B(\R_DATA_TEMPR5[21] ), .C(
        \R_DATA_TEMPR6[21] ), .D(\R_DATA_TEMPR7[21] ), .Y(OR4_973_Y));
    OR4 OR4_806 (.A(OR4_231_Y), .B(OR4_34_Y), .C(OR4_1314_Y), .D(
        OR4_1130_Y), .Y(OR4_806_Y));
    OR4 OR4_701 (.A(OR4_140_Y), .B(OR4_1616_Y), .C(OR4_1001_Y), .D(
        OR4_1530_Y), .Y(OR4_701_Y));
    OR4 \OR4_R_DATA[2]  (.A(OR4_898_Y), .B(OR4_809_Y), .C(OR4_1119_Y), 
        .D(OR4_1242_Y), .Y(R_DATA[2]));
    OR4 OR4_1527 (.A(\R_DATA_TEMPR88[7] ), .B(\R_DATA_TEMPR89[7] ), .C(
        \R_DATA_TEMPR90[7] ), .D(\R_DATA_TEMPR91[7] ), .Y(OR4_1527_Y));
    OR4 OR4_850 (.A(\R_DATA_TEMPR4[12] ), .B(\R_DATA_TEMPR5[12] ), .C(
        \R_DATA_TEMPR6[12] ), .D(\R_DATA_TEMPR7[12] ), .Y(OR4_850_Y));
    OR4 OR4_521 (.A(OR4_1087_Y), .B(OR4_1541_Y), .C(OR4_881_Y), .D(
        OR4_1174_Y), .Y(OR4_521_Y));
    OR4 OR4_1322 (.A(\R_DATA_TEMPR8[26] ), .B(\R_DATA_TEMPR9[26] ), .C(
        \R_DATA_TEMPR10[26] ), .D(\R_DATA_TEMPR11[26] ), .Y(OR4_1322_Y)
        );
    OR4 OR4_876 (.A(\R_DATA_TEMPR56[14] ), .B(\R_DATA_TEMPR57[14] ), 
        .C(\R_DATA_TEMPR58[14] ), .D(\R_DATA_TEMPR59[14] ), .Y(
        OR4_876_Y));
    OR4 OR4_1058 (.A(OR4_742_Y), .B(OR4_555_Y), .C(OR4_183_Y), .D(
        OR4_12_Y), .Y(OR4_1058_Y));
    OR4 OR4_771 (.A(\R_DATA_TEMPR28[32] ), .B(\R_DATA_TEMPR29[32] ), 
        .C(\R_DATA_TEMPR30[32] ), .D(\R_DATA_TEMPR31[32] ), .Y(
        OR4_771_Y));
    OR4 OR4_152 (.A(\R_DATA_TEMPR92[30] ), .B(\R_DATA_TEMPR93[30] ), 
        .C(\R_DATA_TEMPR94[30] ), .D(\R_DATA_TEMPR95[30] ), .Y(
        OR4_152_Y));
    OR4 OR4_893 (.A(\R_DATA_TEMPR16[19] ), .B(\R_DATA_TEMPR17[19] ), 
        .C(\R_DATA_TEMPR18[19] ), .D(\R_DATA_TEMPR19[19] ), .Y(
        OR4_893_Y));
    OR4 OR4_1222 (.A(\R_DATA_TEMPR12[24] ), .B(\R_DATA_TEMPR13[24] ), 
        .C(\R_DATA_TEMPR14[24] ), .D(\R_DATA_TEMPR15[24] ), .Y(
        OR4_1222_Y));
    OR4 OR4_1360 (.A(\R_DATA_TEMPR44[26] ), .B(\R_DATA_TEMPR45[26] ), 
        .C(\R_DATA_TEMPR46[26] ), .D(\R_DATA_TEMPR47[26] ), .Y(
        OR4_1360_Y));
    OR4 OR4_466 (.A(\R_DATA_TEMPR20[11] ), .B(\R_DATA_TEMPR21[11] ), 
        .C(\R_DATA_TEMPR22[11] ), .D(\R_DATA_TEMPR23[11] ), .Y(
        OR4_466_Y));
    OR4 OR4_955 (.A(\R_DATA_TEMPR16[3] ), .B(\R_DATA_TEMPR17[3] ), .C(
        \R_DATA_TEMPR18[3] ), .D(\R_DATA_TEMPR19[3] ), .Y(OR4_955_Y));
    OR4 OR4_39 (.A(\R_DATA_TEMPR24[0] ), .B(\R_DATA_TEMPR25[0] ), .C(
        \R_DATA_TEMPR26[0] ), .D(\R_DATA_TEMPR27[0] ), .Y(OR4_39_Y));
    OR4 OR4_534 (.A(OR4_1613_Y), .B(OR4_290_Y), .C(OR4_1372_Y), .D(
        OR4_593_Y), .Y(OR4_534_Y));
    OR4 OR4_506 (.A(OR4_918_Y), .B(OR4_137_Y), .C(OR4_943_Y), .D(
        OR4_1199_Y), .Y(OR4_506_Y));
    OR4 OR4_211 (.A(\R_DATA_TEMPR12[37] ), .B(\R_DATA_TEMPR13[37] ), 
        .C(\R_DATA_TEMPR14[37] ), .D(\R_DATA_TEMPR15[37] ), .Y(
        OR4_211_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%23%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C0 (.A_DOUT({
        \R_DATA_TEMPR23[39] , \R_DATA_TEMPR23[38] , 
        \R_DATA_TEMPR23[37] , \R_DATA_TEMPR23[36] , 
        \R_DATA_TEMPR23[35] , \R_DATA_TEMPR23[34] , 
        \R_DATA_TEMPR23[33] , \R_DATA_TEMPR23[32] , 
        \R_DATA_TEMPR23[31] , \R_DATA_TEMPR23[30] , 
        \R_DATA_TEMPR23[29] , \R_DATA_TEMPR23[28] , 
        \R_DATA_TEMPR23[27] , \R_DATA_TEMPR23[26] , 
        \R_DATA_TEMPR23[25] , \R_DATA_TEMPR23[24] , 
        \R_DATA_TEMPR23[23] , \R_DATA_TEMPR23[22] , 
        \R_DATA_TEMPR23[21] , \R_DATA_TEMPR23[20] }), .B_DOUT({
        \R_DATA_TEMPR23[19] , \R_DATA_TEMPR23[18] , 
        \R_DATA_TEMPR23[17] , \R_DATA_TEMPR23[16] , 
        \R_DATA_TEMPR23[15] , \R_DATA_TEMPR23[14] , 
        \R_DATA_TEMPR23[13] , \R_DATA_TEMPR23[12] , 
        \R_DATA_TEMPR23[11] , \R_DATA_TEMPR23[10] , 
        \R_DATA_TEMPR23[9] , \R_DATA_TEMPR23[8] , \R_DATA_TEMPR23[7] , 
        \R_DATA_TEMPR23[6] , \R_DATA_TEMPR23[5] , \R_DATA_TEMPR23[4] , 
        \R_DATA_TEMPR23[3] , \R_DATA_TEMPR23[2] , \R_DATA_TEMPR23[1] , 
        \R_DATA_TEMPR23[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1424 (.A(\R_DATA_TEMPR0[3] ), .B(\R_DATA_TEMPR1[3] ), .C(
        \R_DATA_TEMPR2[3] ), .D(\R_DATA_TEMPR3[3] ), .Y(OR4_1424_Y));
    OR4 OR4_932 (.A(\R_DATA_TEMPR0[39] ), .B(\R_DATA_TEMPR1[39] ), .C(
        \R_DATA_TEMPR2[39] ), .D(\R_DATA_TEMPR3[39] ), .Y(OR4_932_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%2%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C0 (.A_DOUT({
        \R_DATA_TEMPR2[39] , \R_DATA_TEMPR2[38] , \R_DATA_TEMPR2[37] , 
        \R_DATA_TEMPR2[36] , \R_DATA_TEMPR2[35] , \R_DATA_TEMPR2[34] , 
        \R_DATA_TEMPR2[33] , \R_DATA_TEMPR2[32] , \R_DATA_TEMPR2[31] , 
        \R_DATA_TEMPR2[30] , \R_DATA_TEMPR2[29] , \R_DATA_TEMPR2[28] , 
        \R_DATA_TEMPR2[27] , \R_DATA_TEMPR2[26] , \R_DATA_TEMPR2[25] , 
        \R_DATA_TEMPR2[24] , \R_DATA_TEMPR2[23] , \R_DATA_TEMPR2[22] , 
        \R_DATA_TEMPR2[21] , \R_DATA_TEMPR2[20] }), .B_DOUT({
        \R_DATA_TEMPR2[19] , \R_DATA_TEMPR2[18] , \R_DATA_TEMPR2[17] , 
        \R_DATA_TEMPR2[16] , \R_DATA_TEMPR2[15] , \R_DATA_TEMPR2[14] , 
        \R_DATA_TEMPR2[13] , \R_DATA_TEMPR2[12] , \R_DATA_TEMPR2[11] , 
        \R_DATA_TEMPR2[10] , \R_DATA_TEMPR2[9] , \R_DATA_TEMPR2[8] , 
        \R_DATA_TEMPR2[7] , \R_DATA_TEMPR2[6] , \R_DATA_TEMPR2[5] , 
        \R_DATA_TEMPR2[4] , \R_DATA_TEMPR2[3] , \R_DATA_TEMPR2[2] , 
        \R_DATA_TEMPR2[1] , \R_DATA_TEMPR2[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[2][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR2 OR2_9 (.A(\R_DATA_TEMPR84[24] ), .B(\R_DATA_TEMPR85[24] ), .Y(
        OR2_9_Y));
    OR4 OR4_484 (.A(\R_DATA_TEMPR48[20] ), .B(\R_DATA_TEMPR49[20] ), 
        .C(\R_DATA_TEMPR50[20] ), .D(\R_DATA_TEMPR51[20] ), .Y(
        OR4_484_Y));
    OR4 OR4_1552 (.A(\R_DATA_TEMPR112[26] ), .B(\R_DATA_TEMPR113[26] ), 
        .C(\R_DATA_TEMPR114[26] ), .D(\R_DATA_TEMPR115[26] ), .Y(
        OR4_1552_Y));
    OR4 OR4_1014 (.A(\R_DATA_TEMPR4[33] ), .B(\R_DATA_TEMPR5[33] ), .C(
        \R_DATA_TEMPR6[33] ), .D(\R_DATA_TEMPR7[33] ), .Y(OR4_1014_Y));
    OR4 OR4_1435 (.A(OR4_436_Y), .B(OR4_1387_Y), .C(OR4_1463_Y), .D(
        OR4_646_Y), .Y(OR4_1435_Y));
    OR4 OR4_1190 (.A(\R_DATA_TEMPR20[33] ), .B(\R_DATA_TEMPR21[33] ), 
        .C(\R_DATA_TEMPR22[33] ), .D(\R_DATA_TEMPR23[33] ), .Y(
        OR4_1190_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%120%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R120C0 (.A_DOUT({
        \R_DATA_TEMPR120[39] , \R_DATA_TEMPR120[38] , 
        \R_DATA_TEMPR120[37] , \R_DATA_TEMPR120[36] , 
        \R_DATA_TEMPR120[35] , \R_DATA_TEMPR120[34] , 
        \R_DATA_TEMPR120[33] , \R_DATA_TEMPR120[32] , 
        \R_DATA_TEMPR120[31] , \R_DATA_TEMPR120[30] , 
        \R_DATA_TEMPR120[29] , \R_DATA_TEMPR120[28] , 
        \R_DATA_TEMPR120[27] , \R_DATA_TEMPR120[26] , 
        \R_DATA_TEMPR120[25] , \R_DATA_TEMPR120[24] , 
        \R_DATA_TEMPR120[23] , \R_DATA_TEMPR120[22] , 
        \R_DATA_TEMPR120[21] , \R_DATA_TEMPR120[20] }), .B_DOUT({
        \R_DATA_TEMPR120[19] , \R_DATA_TEMPR120[18] , 
        \R_DATA_TEMPR120[17] , \R_DATA_TEMPR120[16] , 
        \R_DATA_TEMPR120[15] , \R_DATA_TEMPR120[14] , 
        \R_DATA_TEMPR120[13] , \R_DATA_TEMPR120[12] , 
        \R_DATA_TEMPR120[11] , \R_DATA_TEMPR120[10] , 
        \R_DATA_TEMPR120[9] , \R_DATA_TEMPR120[8] , 
        \R_DATA_TEMPR120[7] , \R_DATA_TEMPR120[6] , 
        \R_DATA_TEMPR120[5] , \R_DATA_TEMPR120[4] , 
        \R_DATA_TEMPR120[3] , \R_DATA_TEMPR120[2] , 
        \R_DATA_TEMPR120[1] , \R_DATA_TEMPR120[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[120][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[30] , \BLKY1[0] , \BLKY0[0] }), 
        .A_CLK(CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], 
        W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], 
        W_DATA[31], W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], 
        W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], 
        W_DATA[21], W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], 
        WBYTE_EN[2]}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], 
        W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], 
        W_ADDR[0], GND, GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[30] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA[19], 
        W_DATA[18], W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], 
        W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], W_DATA[9], 
        W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], 
        W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_576 (.A(OR4_1568_Y), .B(OR4_383_Y), .C(OR4_364_Y), .D(
        OR4_1125_Y), .Y(OR4_576_Y));
    OR4 OR4_1470 (.A(OR4_124_Y), .B(OR4_1269_Y), .C(OR4_1330_Y), .D(
        OR4_721_Y), .Y(OR4_1470_Y));
    OR4 OR4_1224 (.A(\R_DATA_TEMPR40[25] ), .B(\R_DATA_TEMPR41[25] ), 
        .C(\R_DATA_TEMPR42[25] ), .D(\R_DATA_TEMPR43[25] ), .Y(
        OR4_1224_Y));
    OR4 OR4_145 (.A(\R_DATA_TEMPR104[26] ), .B(\R_DATA_TEMPR105[26] ), 
        .C(\R_DATA_TEMPR106[26] ), .D(\R_DATA_TEMPR107[26] ), .Y(
        OR4_145_Y));
    OR4 OR4_362 (.A(\R_DATA_TEMPR92[7] ), .B(\R_DATA_TEMPR93[7] ), .C(
        \R_DATA_TEMPR94[7] ), .D(\R_DATA_TEMPR95[7] ), .Y(OR4_362_Y));
    OR4 OR4_222 (.A(\R_DATA_TEMPR68[38] ), .B(\R_DATA_TEMPR69[38] ), 
        .C(\R_DATA_TEMPR70[38] ), .D(\R_DATA_TEMPR71[38] ), .Y(
        OR4_222_Y));
    OR4 OR4_1313 (.A(\R_DATA_TEMPR76[20] ), .B(\R_DATA_TEMPR77[20] ), 
        .C(\R_DATA_TEMPR78[20] ), .D(\R_DATA_TEMPR79[20] ), .Y(
        OR4_1313_Y));
    OR4 OR4_1143 (.A(\R_DATA_TEMPR0[27] ), .B(\R_DATA_TEMPR1[27] ), .C(
        \R_DATA_TEMPR2[27] ), .D(\R_DATA_TEMPR3[27] ), .Y(OR4_1143_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%32%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R32C0 (.A_DOUT({
        \R_DATA_TEMPR32[39] , \R_DATA_TEMPR32[38] , 
        \R_DATA_TEMPR32[37] , \R_DATA_TEMPR32[36] , 
        \R_DATA_TEMPR32[35] , \R_DATA_TEMPR32[34] , 
        \R_DATA_TEMPR32[33] , \R_DATA_TEMPR32[32] , 
        \R_DATA_TEMPR32[31] , \R_DATA_TEMPR32[30] , 
        \R_DATA_TEMPR32[29] , \R_DATA_TEMPR32[28] , 
        \R_DATA_TEMPR32[27] , \R_DATA_TEMPR32[26] , 
        \R_DATA_TEMPR32[25] , \R_DATA_TEMPR32[24] , 
        \R_DATA_TEMPR32[23] , \R_DATA_TEMPR32[22] , 
        \R_DATA_TEMPR32[21] , \R_DATA_TEMPR32[20] }), .B_DOUT({
        \R_DATA_TEMPR32[19] , \R_DATA_TEMPR32[18] , 
        \R_DATA_TEMPR32[17] , \R_DATA_TEMPR32[16] , 
        \R_DATA_TEMPR32[15] , \R_DATA_TEMPR32[14] , 
        \R_DATA_TEMPR32[13] , \R_DATA_TEMPR32[12] , 
        \R_DATA_TEMPR32[11] , \R_DATA_TEMPR32[10] , 
        \R_DATA_TEMPR32[9] , \R_DATA_TEMPR32[8] , \R_DATA_TEMPR32[7] , 
        \R_DATA_TEMPR32[6] , \R_DATA_TEMPR32[5] , \R_DATA_TEMPR32[4] , 
        \R_DATA_TEMPR32[3] , \R_DATA_TEMPR32[2] , \R_DATA_TEMPR32[1] , 
        \R_DATA_TEMPR32[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[32][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[8] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[8] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_16 (.A(\R_DATA_TEMPR104[34] ), .B(\R_DATA_TEMPR105[34] ), 
        .C(\R_DATA_TEMPR106[34] ), .D(\R_DATA_TEMPR107[34] ), .Y(
        OR4_16_Y));
    OR4 OR4_386 (.A(OR4_1260_Y), .B(OR4_512_Y), .C(OR4_480_Y), .D(
        OR4_1256_Y), .Y(OR4_386_Y));
    OR4 OR4_1327 (.A(OR4_549_Y), .B(OR2_5_Y), .C(\R_DATA_TEMPR86[39] ), 
        .D(\R_DATA_TEMPR87[39] ), .Y(OR4_1327_Y));
    OR4 OR4_447 (.A(\R_DATA_TEMPR68[27] ), .B(\R_DATA_TEMPR69[27] ), 
        .C(\R_DATA_TEMPR70[27] ), .D(\R_DATA_TEMPR71[27] ), .Y(
        OR4_447_Y));
    OR4 OR4_259 (.A(\R_DATA_TEMPR8[1] ), .B(\R_DATA_TEMPR9[1] ), .C(
        \R_DATA_TEMPR10[1] ), .D(\R_DATA_TEMPR11[1] ), .Y(OR4_259_Y));
    OR4 OR4_4 (.A(\R_DATA_TEMPR96[27] ), .B(\R_DATA_TEMPR97[27] ), .C(
        \R_DATA_TEMPR98[27] ), .D(\R_DATA_TEMPR99[27] ), .Y(OR4_4_Y));
    OR4 OR4_331 (.A(\R_DATA_TEMPR32[20] ), .B(\R_DATA_TEMPR33[20] ), 
        .C(\R_DATA_TEMPR34[20] ), .D(\R_DATA_TEMPR35[20] ), .Y(
        OR4_331_Y));
    OR4 OR4_1605 (.A(\R_DATA_TEMPR16[23] ), .B(\R_DATA_TEMPR17[23] ), 
        .C(\R_DATA_TEMPR18[23] ), .D(\R_DATA_TEMPR19[23] ), .Y(
        OR4_1605_Y));
    OR4 OR4_1171 (.A(OR4_1491_Y), .B(OR4_806_Y), .C(OR4_1138_Y), .D(
        OR4_345_Y), .Y(OR4_1171_Y));
    OR4 OR4_512 (.A(\R_DATA_TEMPR36[17] ), .B(\R_DATA_TEMPR37[17] ), 
        .C(\R_DATA_TEMPR38[17] ), .D(\R_DATA_TEMPR39[17] ), .Y(
        OR4_512_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%77%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R77C0 (.A_DOUT({
        \R_DATA_TEMPR77[39] , \R_DATA_TEMPR77[38] , 
        \R_DATA_TEMPR77[37] , \R_DATA_TEMPR77[36] , 
        \R_DATA_TEMPR77[35] , \R_DATA_TEMPR77[34] , 
        \R_DATA_TEMPR77[33] , \R_DATA_TEMPR77[32] , 
        \R_DATA_TEMPR77[31] , \R_DATA_TEMPR77[30] , 
        \R_DATA_TEMPR77[29] , \R_DATA_TEMPR77[28] , 
        \R_DATA_TEMPR77[27] , \R_DATA_TEMPR77[26] , 
        \R_DATA_TEMPR77[25] , \R_DATA_TEMPR77[24] , 
        \R_DATA_TEMPR77[23] , \R_DATA_TEMPR77[22] , 
        \R_DATA_TEMPR77[21] , \R_DATA_TEMPR77[20] }), .B_DOUT({
        \R_DATA_TEMPR77[19] , \R_DATA_TEMPR77[18] , 
        \R_DATA_TEMPR77[17] , \R_DATA_TEMPR77[16] , 
        \R_DATA_TEMPR77[15] , \R_DATA_TEMPR77[14] , 
        \R_DATA_TEMPR77[13] , \R_DATA_TEMPR77[12] , 
        \R_DATA_TEMPR77[11] , \R_DATA_TEMPR77[10] , 
        \R_DATA_TEMPR77[9] , \R_DATA_TEMPR77[8] , \R_DATA_TEMPR77[7] , 
        \R_DATA_TEMPR77[6] , \R_DATA_TEMPR77[5] , \R_DATA_TEMPR77[4] , 
        \R_DATA_TEMPR77[3] , \R_DATA_TEMPR77[2] , \R_DATA_TEMPR77[1] , 
        \R_DATA_TEMPR77[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[77][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[19] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[19] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1549 (.A(OR4_581_Y), .B(OR4_1363_Y), .C(OR4_185_Y), .D(
        OR4_507_Y), .Y(OR4_1549_Y));
    OR4 OR4_1207 (.A(\R_DATA_TEMPR20[21] ), .B(\R_DATA_TEMPR21[21] ), 
        .C(\R_DATA_TEMPR22[21] ), .D(\R_DATA_TEMPR23[21] ), .Y(
        OR4_1207_Y));
    OR4 OR4_320 (.A(\R_DATA_TEMPR44[18] ), .B(\R_DATA_TEMPR45[18] ), 
        .C(\R_DATA_TEMPR46[18] ), .D(\R_DATA_TEMPR47[18] ), .Y(
        OR4_320_Y));
    OR4 OR4_1576 (.A(\R_DATA_TEMPR88[24] ), .B(\R_DATA_TEMPR89[24] ), 
        .C(\R_DATA_TEMPR90[24] ), .D(\R_DATA_TEMPR91[24] ), .Y(
        OR4_1576_Y));
    OR4 OR4_430 (.A(OR4_1422_Y), .B(OR2_6_Y), .C(\R_DATA_TEMPR86[3] ), 
        .D(\R_DATA_TEMPR87[3] ), .Y(OR4_430_Y));
    OR4 OR4_1634 (.A(\R_DATA_TEMPR80[34] ), .B(\R_DATA_TEMPR81[34] ), 
        .C(\R_DATA_TEMPR82[34] ), .D(\R_DATA_TEMPR83[34] ), .Y(
        OR4_1634_Y));
    OR4 OR4_1265 (.A(\R_DATA_TEMPR92[18] ), .B(\R_DATA_TEMPR93[18] ), 
        .C(\R_DATA_TEMPR94[18] ), .D(\R_DATA_TEMPR95[18] ), .Y(
        OR4_1265_Y));
    OR4 \OR4_R_DATA[14]  (.A(OR4_1551_Y), .B(OR4_979_Y), .C(OR4_135_Y), 
        .D(OR4_861_Y), .Y(R_DATA[14]));
    OR4 OR4_595 (.A(\R_DATA_TEMPR72[32] ), .B(\R_DATA_TEMPR73[32] ), 
        .C(\R_DATA_TEMPR74[32] ), .D(\R_DATA_TEMPR75[32] ), .Y(
        OR4_595_Y));
    OR4 OR4_245 (.A(\R_DATA_TEMPR24[10] ), .B(\R_DATA_TEMPR25[10] ), 
        .C(\R_DATA_TEMPR26[10] ), .D(\R_DATA_TEMPR27[10] ), .Y(
        OR4_245_Y));
    OR4 OR4_508 (.A(OR4_958_Y), .B(OR2_18_Y), .C(\R_DATA_TEMPR86[30] ), 
        .D(\R_DATA_TEMPR87[30] ), .Y(OR4_508_Y));
    OR4 OR4_1561 (.A(OR4_1153_Y), .B(OR2_24_Y), .C(
        \R_DATA_TEMPR86[36] ), .D(\R_DATA_TEMPR87[36] ), .Y(OR4_1561_Y)
        );
    OR4 OR4_1390 (.A(\R_DATA_TEMPR32[27] ), .B(\R_DATA_TEMPR33[27] ), 
        .C(\R_DATA_TEMPR34[27] ), .D(\R_DATA_TEMPR35[27] ), .Y(
        OR4_1390_Y));
    OR4 OR4_50 (.A(\R_DATA_TEMPR124[25] ), .B(\R_DATA_TEMPR125[25] ), 
        .C(\R_DATA_TEMPR126[25] ), .D(\R_DATA_TEMPR127[25] ), .Y(
        OR4_50_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%87%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R87C0 (.A_DOUT({
        \R_DATA_TEMPR87[39] , \R_DATA_TEMPR87[38] , 
        \R_DATA_TEMPR87[37] , \R_DATA_TEMPR87[36] , 
        \R_DATA_TEMPR87[35] , \R_DATA_TEMPR87[34] , 
        \R_DATA_TEMPR87[33] , \R_DATA_TEMPR87[32] , 
        \R_DATA_TEMPR87[31] , \R_DATA_TEMPR87[30] , 
        \R_DATA_TEMPR87[29] , \R_DATA_TEMPR87[28] , 
        \R_DATA_TEMPR87[27] , \R_DATA_TEMPR87[26] , 
        \R_DATA_TEMPR87[25] , \R_DATA_TEMPR87[24] , 
        \R_DATA_TEMPR87[23] , \R_DATA_TEMPR87[22] , 
        \R_DATA_TEMPR87[21] , \R_DATA_TEMPR87[20] }), .B_DOUT({
        \R_DATA_TEMPR87[19] , \R_DATA_TEMPR87[18] , 
        \R_DATA_TEMPR87[17] , \R_DATA_TEMPR87[16] , 
        \R_DATA_TEMPR87[15] , \R_DATA_TEMPR87[14] , 
        \R_DATA_TEMPR87[13] , \R_DATA_TEMPR87[12] , 
        \R_DATA_TEMPR87[11] , \R_DATA_TEMPR87[10] , 
        \R_DATA_TEMPR87[9] , \R_DATA_TEMPR87[8] , \R_DATA_TEMPR87[7] , 
        \R_DATA_TEMPR87[6] , \R_DATA_TEMPR87[5] , \R_DATA_TEMPR87[4] , 
        \R_DATA_TEMPR87[3] , \R_DATA_TEMPR87[2] , \R_DATA_TEMPR87[1] , 
        \R_DATA_TEMPR87[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[87][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[21] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[21] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1602 (.A(\R_DATA_TEMPR96[15] ), .B(\R_DATA_TEMPR97[15] ), 
        .C(\R_DATA_TEMPR98[15] ), .D(\R_DATA_TEMPR99[15] ), .Y(
        OR4_1602_Y));
    OR4 OR4_842 (.A(\R_DATA_TEMPR76[7] ), .B(\R_DATA_TEMPR77[7] ), .C(
        \R_DATA_TEMPR78[7] ), .D(\R_DATA_TEMPR79[7] ), .Y(OR4_842_Y));
    OR4 OR4_1406 (.A(\R_DATA_TEMPR48[33] ), .B(\R_DATA_TEMPR49[33] ), 
        .C(\R_DATA_TEMPR50[33] ), .D(\R_DATA_TEMPR51[33] ), .Y(
        OR4_1406_Y));
    OR4 OR4_1304 (.A(\R_DATA_TEMPR24[6] ), .B(\R_DATA_TEMPR25[6] ), .C(
        \R_DATA_TEMPR26[6] ), .D(\R_DATA_TEMPR27[6] ), .Y(OR4_1304_Y));
    OR4 OR4_859 (.A(\R_DATA_TEMPR60[25] ), .B(\R_DATA_TEMPR61[25] ), 
        .C(\R_DATA_TEMPR62[25] ), .D(\R_DATA_TEMPR63[25] ), .Y(
        OR4_859_Y));
    OR4 OR4_823 (.A(\R_DATA_TEMPR40[39] ), .B(\R_DATA_TEMPR41[39] ), 
        .C(\R_DATA_TEMPR42[39] ), .D(\R_DATA_TEMPR43[39] ), .Y(
        OR4_823_Y));
    OR4 OR4_514 (.A(\R_DATA_TEMPR44[39] ), .B(\R_DATA_TEMPR45[39] ), 
        .C(\R_DATA_TEMPR46[39] ), .D(\R_DATA_TEMPR47[39] ), .Y(
        OR4_514_Y));
    OR4 OR4_1336 (.A(\R_DATA_TEMPR72[15] ), .B(\R_DATA_TEMPR73[15] ), 
        .C(\R_DATA_TEMPR74[15] ), .D(\R_DATA_TEMPR75[15] ), .Y(
        OR4_1336_Y));
    OR4 OR4_578 (.A(\R_DATA_TEMPR28[15] ), .B(\R_DATA_TEMPR29[15] ), 
        .C(\R_DATA_TEMPR30[15] ), .D(\R_DATA_TEMPR31[15] ), .Y(
        OR4_578_Y));
    OR4 OR4_693 (.A(\R_DATA_TEMPR88[38] ), .B(\R_DATA_TEMPR89[38] ), 
        .C(\R_DATA_TEMPR90[38] ), .D(\R_DATA_TEMPR91[38] ), .Y(
        OR4_693_Y));
    OR4 OR4_57 (.A(\R_DATA_TEMPR32[11] ), .B(\R_DATA_TEMPR33[11] ), .C(
        \R_DATA_TEMPR34[11] ), .D(\R_DATA_TEMPR35[11] ), .Y(OR4_57_Y));
    OR4 OR4_32 (.A(\R_DATA_TEMPR100[12] ), .B(\R_DATA_TEMPR101[12] ), 
        .C(\R_DATA_TEMPR102[12] ), .D(\R_DATA_TEMPR103[12] ), .Y(
        OR4_32_Y));
    OR4 OR4_260 (.A(\R_DATA_TEMPR48[28] ), .B(\R_DATA_TEMPR49[28] ), 
        .C(\R_DATA_TEMPR50[28] ), .D(\R_DATA_TEMPR51[28] ), .Y(
        OR4_260_Y));
    OR4 OR4_912 (.A(\R_DATA_TEMPR44[15] ), .B(\R_DATA_TEMPR45[15] ), 
        .C(\R_DATA_TEMPR46[15] ), .D(\R_DATA_TEMPR47[15] ), .Y(
        OR4_912_Y));
    OR4 OR4_567 (.A(\R_DATA_TEMPR12[1] ), .B(\R_DATA_TEMPR13[1] ), .C(
        \R_DATA_TEMPR14[1] ), .D(\R_DATA_TEMPR15[1] ), .Y(OR4_567_Y));
    OR4 OR4_1631 (.A(\R_DATA_TEMPR24[7] ), .B(\R_DATA_TEMPR25[7] ), .C(
        \R_DATA_TEMPR26[7] ), .D(\R_DATA_TEMPR27[7] ), .Y(OR4_1631_Y));
    OR4 OR4_1477 (.A(\R_DATA_TEMPR88[2] ), .B(\R_DATA_TEMPR89[2] ), .C(
        \R_DATA_TEMPR90[2] ), .D(\R_DATA_TEMPR91[2] ), .Y(OR4_1477_Y));
    OR4 OR4_1057 (.A(\R_DATA_TEMPR4[26] ), .B(\R_DATA_TEMPR5[26] ), .C(
        \R_DATA_TEMPR6[26] ), .D(\R_DATA_TEMPR7[26] ), .Y(OR4_1057_Y));
    OR4 OR4_1425 (.A(OR4_37_Y), .B(OR4_1057_Y), .C(OR4_1322_Y), .D(
        OR4_263_Y), .Y(OR4_1425_Y));
    OR4 OR4_1287 (.A(OR4_1281_Y), .B(OR2_1_Y), .C(\R_DATA_TEMPR86[4] ), 
        .D(\R_DATA_TEMPR87[4] ), .Y(OR4_1287_Y));
    OR4 OR4_1607 (.A(\R_DATA_TEMPR48[26] ), .B(\R_DATA_TEMPR49[26] ), 
        .C(\R_DATA_TEMPR50[26] ), .D(\R_DATA_TEMPR51[26] ), .Y(
        OR4_1607_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%122%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R122C0 (.A_DOUT({
        \R_DATA_TEMPR122[39] , \R_DATA_TEMPR122[38] , 
        \R_DATA_TEMPR122[37] , \R_DATA_TEMPR122[36] , 
        \R_DATA_TEMPR122[35] , \R_DATA_TEMPR122[34] , 
        \R_DATA_TEMPR122[33] , \R_DATA_TEMPR122[32] , 
        \R_DATA_TEMPR122[31] , \R_DATA_TEMPR122[30] , 
        \R_DATA_TEMPR122[29] , \R_DATA_TEMPR122[28] , 
        \R_DATA_TEMPR122[27] , \R_DATA_TEMPR122[26] , 
        \R_DATA_TEMPR122[25] , \R_DATA_TEMPR122[24] , 
        \R_DATA_TEMPR122[23] , \R_DATA_TEMPR122[22] , 
        \R_DATA_TEMPR122[21] , \R_DATA_TEMPR122[20] }), .B_DOUT({
        \R_DATA_TEMPR122[19] , \R_DATA_TEMPR122[18] , 
        \R_DATA_TEMPR122[17] , \R_DATA_TEMPR122[16] , 
        \R_DATA_TEMPR122[15] , \R_DATA_TEMPR122[14] , 
        \R_DATA_TEMPR122[13] , \R_DATA_TEMPR122[12] , 
        \R_DATA_TEMPR122[11] , \R_DATA_TEMPR122[10] , 
        \R_DATA_TEMPR122[9] , \R_DATA_TEMPR122[8] , 
        \R_DATA_TEMPR122[7] , \R_DATA_TEMPR122[6] , 
        \R_DATA_TEMPR122[5] , \R_DATA_TEMPR122[4] , 
        \R_DATA_TEMPR122[3] , \R_DATA_TEMPR122[2] , 
        \R_DATA_TEMPR122[1] , \R_DATA_TEMPR122[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[122][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[30] , R_ADDR[10], \BLKY0[0] }), 
        .A_CLK(CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], 
        W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], 
        W_DATA[31], W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], 
        W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], 
        W_DATA[21], W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], 
        WBYTE_EN[2]}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], 
        W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], 
        W_ADDR[0], GND, GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[30] , 
        W_ADDR[10], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA[19], 
        W_DATA[18], W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], 
        W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], W_DATA[9], 
        W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], 
        W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_406 (.A(\R_DATA_TEMPR52[17] ), .B(\R_DATA_TEMPR53[17] ), 
        .C(\R_DATA_TEMPR54[17] ), .D(\R_DATA_TEMPR55[17] ), .Y(
        OR4_406_Y));
    OR4 OR4_1016 (.A(OR4_78_Y), .B(OR4_387_Y), .C(OR4_1476_Y), .D(
        OR4_682_Y), .Y(OR4_1016_Y));
    OR4 OR4_1630 (.A(\R_DATA_TEMPR108[33] ), .B(\R_DATA_TEMPR109[33] ), 
        .C(\R_DATA_TEMPR110[33] ), .D(\R_DATA_TEMPR111[33] ), .Y(
        OR4_1630_Y));
    OR4 OR4_1075 (.A(OR4_740_Y), .B(OR4_990_Y), .C(OR4_1177_Y), .D(
        OR4_1255_Y), .Y(OR4_1075_Y));
    OR4 OR4_443 (.A(\R_DATA_TEMPR52[11] ), .B(\R_DATA_TEMPR53[11] ), 
        .C(\R_DATA_TEMPR54[11] ), .D(\R_DATA_TEMPR55[11] ), .Y(
        OR4_443_Y));
    OR4 OR4_669 (.A(\R_DATA_TEMPR60[39] ), .B(\R_DATA_TEMPR61[39] ), 
        .C(\R_DATA_TEMPR62[39] ), .D(\R_DATA_TEMPR63[39] ), .Y(
        OR4_669_Y));
    OR4 OR4_641 (.A(\R_DATA_TEMPR56[17] ), .B(\R_DATA_TEMPR57[17] ), 
        .C(\R_DATA_TEMPR58[17] ), .D(\R_DATA_TEMPR59[17] ), .Y(
        OR4_641_Y));
    OR4 OR4_184 (.A(\R_DATA_TEMPR0[29] ), .B(\R_DATA_TEMPR1[29] ), .C(
        \R_DATA_TEMPR2[29] ), .D(\R_DATA_TEMPR3[29] ), .Y(OR4_184_Y));
    OR4 OR4_311 (.A(OR4_598_Y), .B(OR4_1623_Y), .C(OR4_235_Y), .D(
        OR4_804_Y), .Y(OR4_311_Y));
    OR4 OR4_476 (.A(\R_DATA_TEMPR92[16] ), .B(\R_DATA_TEMPR93[16] ), 
        .C(\R_DATA_TEMPR94[16] ), .D(\R_DATA_TEMPR95[16] ), .Y(
        OR4_476_Y));
    OR4 OR4_248 (.A(OR4_418_Y), .B(OR2_35_Y), .C(\R_DATA_TEMPR86[26] ), 
        .D(\R_DATA_TEMPR87[26] ), .Y(OR4_248_Y));
    OR4 OR4_1486 (.A(\R_DATA_TEMPR48[38] ), .B(\R_DATA_TEMPR49[38] ), 
        .C(\R_DATA_TEMPR50[38] ), .D(\R_DATA_TEMPR51[38] ), .Y(
        OR4_1486_Y));
    OR4 OR4_1384 (.A(\R_DATA_TEMPR104[27] ), .B(\R_DATA_TEMPR105[27] ), 
        .C(\R_DATA_TEMPR106[27] ), .D(\R_DATA_TEMPR107[27] ), .Y(
        OR4_1384_Y));
    OR4 OR4_999 (.A(\R_DATA_TEMPR104[2] ), .B(\R_DATA_TEMPR105[2] ), 
        .C(\R_DATA_TEMPR106[2] ), .D(\R_DATA_TEMPR107[2] ), .Y(
        OR4_999_Y));
    OR4 OR4_990 (.A(\R_DATA_TEMPR68[8] ), .B(\R_DATA_TEMPR69[8] ), .C(
        \R_DATA_TEMPR70[8] ), .D(\R_DATA_TEMPR71[8] ), .Y(OR4_990_Y));
    OR4 OR4_1311 (.A(\R_DATA_TEMPR48[9] ), .B(\R_DATA_TEMPR49[9] ), .C(
        \R_DATA_TEMPR50[9] ), .D(\R_DATA_TEMPR51[9] ), .Y(OR4_1311_Y));
    OR4 OR4_757 (.A(OR4_1278_Y), .B(OR4_509_Y), .C(OR4_1304_Y), .D(
        OR4_1556_Y), .Y(OR4_757_Y));
    OR4 OR4_1309 (.A(\R_DATA_TEMPR80[15] ), .B(\R_DATA_TEMPR81[15] ), 
        .C(\R_DATA_TEMPR82[15] ), .D(\R_DATA_TEMPR83[15] ), .Y(
        OR4_1309_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[30]  (.A(CFG3_1_Y), .B(CFG3_3_Y)
        , .Y(\BLKY2[30] ));
    OR4 OR4_754 (.A(\R_DATA_TEMPR36[3] ), .B(\R_DATA_TEMPR37[3] ), .C(
        \R_DATA_TEMPR38[3] ), .D(\R_DATA_TEMPR39[3] ), .Y(OR4_754_Y));
    OR4 OR4_302 (.A(\R_DATA_TEMPR108[7] ), .B(\R_DATA_TEMPR109[7] ), 
        .C(\R_DATA_TEMPR110[7] ), .D(\R_DATA_TEMPR111[7] ), .Y(
        OR4_302_Y));
    OR4 OR4_266 (.A(\R_DATA_TEMPR32[26] ), .B(\R_DATA_TEMPR33[26] ), 
        .C(\R_DATA_TEMPR34[26] ), .D(\R_DATA_TEMPR35[26] ), .Y(
        OR4_266_Y));
    OR4 OR4_1545 (.A(\R_DATA_TEMPR44[4] ), .B(\R_DATA_TEMPR45[4] ), .C(
        \R_DATA_TEMPR46[4] ), .D(\R_DATA_TEMPR47[4] ), .Y(OR4_1545_Y));
    OR4 OR4_1295 (.A(\R_DATA_TEMPR88[39] ), .B(\R_DATA_TEMPR89[39] ), 
        .C(\R_DATA_TEMPR90[39] ), .D(\R_DATA_TEMPR91[39] ), .Y(
        OR4_1295_Y));
    OR4 OR4_1000 (.A(\R_DATA_TEMPR120[26] ), .B(\R_DATA_TEMPR121[26] ), 
        .C(\R_DATA_TEMPR122[26] ), .D(\R_DATA_TEMPR123[26] ), .Y(
        OR4_1000_Y));
    OR4 OR4_10 (.A(OR4_403_Y), .B(OR4_1359_Y), .C(OR4_1332_Y), .D(
        OR4_476_Y), .Y(OR4_10_Y));
    OR4 OR4_25 (.A(\R_DATA_TEMPR28[27] ), .B(\R_DATA_TEMPR29[27] ), .C(
        \R_DATA_TEMPR30[27] ), .D(\R_DATA_TEMPR31[27] ), .Y(OR4_25_Y));
    OR4 OR4_76 (.A(\R_DATA_TEMPR52[5] ), .B(\R_DATA_TEMPR53[5] ), .C(
        \R_DATA_TEMPR54[5] ), .D(\R_DATA_TEMPR55[5] ), .Y(OR4_76_Y));
    OR4 OR4_410 (.A(OR4_116_Y), .B(OR4_1592_Y), .C(OR4_87_Y), .D(
        OR4_35_Y), .Y(OR4_410_Y));
    OR4 OR4_1624 (.A(\R_DATA_TEMPR4[23] ), .B(\R_DATA_TEMPR5[23] ), .C(
        \R_DATA_TEMPR6[23] ), .D(\R_DATA_TEMPR7[23] ), .Y(OR4_1624_Y));
    OR4 OR4_983 (.A(\R_DATA_TEMPR48[10] ), .B(\R_DATA_TEMPR49[10] ), 
        .C(\R_DATA_TEMPR50[10] ), .D(\R_DATA_TEMPR51[10] ), .Y(
        OR4_983_Y));
    OR4 OR4_339 (.A(\R_DATA_TEMPR88[32] ), .B(\R_DATA_TEMPR89[32] ), 
        .C(\R_DATA_TEMPR90[32] ), .D(\R_DATA_TEMPR91[32] ), .Y(
        OR4_339_Y));
    OR4 OR4_193 (.A(\R_DATA_TEMPR72[33] ), .B(\R_DATA_TEMPR73[33] ), 
        .C(\R_DATA_TEMPR74[33] ), .D(\R_DATA_TEMPR75[33] ), .Y(
        OR4_193_Y));
    OR4 OR4_1591 (.A(OR4_668_Y), .B(OR4_1190_Y), .C(OR4_695_Y), .D(
        OR4_206_Y), .Y(OR4_1591_Y));
    OR4 OR4_1438 (.A(\R_DATA_TEMPR116[15] ), .B(\R_DATA_TEMPR117[15] ), 
        .C(\R_DATA_TEMPR118[15] ), .D(\R_DATA_TEMPR119[15] ), .Y(
        OR4_1438_Y));
    OR4 OR4_372 (.A(\R_DATA_TEMPR36[35] ), .B(\R_DATA_TEMPR37[35] ), 
        .C(\R_DATA_TEMPR38[35] ), .D(\R_DATA_TEMPR39[35] ), .Y(
        OR4_372_Y));
    OR4 OR4_1246 (.A(\R_DATA_TEMPR92[9] ), .B(\R_DATA_TEMPR93[9] ), .C(
        \R_DATA_TEMPR94[9] ), .D(\R_DATA_TEMPR95[9] ), .Y(OR4_1246_Y));
    OR4 OR4_851 (.A(OR4_1282_Y), .B(OR4_1025_Y), .C(OR4_1576_Y), .D(
        OR4_969_Y), .Y(OR4_851_Y));
    OR4 OR4_525 (.A(\R_DATA_TEMPR124[11] ), .B(\R_DATA_TEMPR125[11] ), 
        .C(\R_DATA_TEMPR126[11] ), .D(\R_DATA_TEMPR127[11] ), .Y(
        OR4_525_Y));
    OR4 OR4_17 (.A(\R_DATA_TEMPR72[1] ), .B(\R_DATA_TEMPR73[1] ), .C(
        \R_DATA_TEMPR74[1] ), .D(\R_DATA_TEMPR75[1] ), .Y(OR4_17_Y));
    OR4 OR4_886 (.A(\R_DATA_TEMPR48[4] ), .B(\R_DATA_TEMPR49[4] ), .C(
        \R_DATA_TEMPR50[4] ), .D(\R_DATA_TEMPR51[4] ), .Y(OR4_886_Y));
    OR4 OR4_781 (.A(\R_DATA_TEMPR116[3] ), .B(\R_DATA_TEMPR117[3] ), 
        .C(\R_DATA_TEMPR118[3] ), .D(\R_DATA_TEMPR119[3] ), .Y(
        OR4_781_Y));
    OR4 OR4_664 (.A(\R_DATA_TEMPR124[10] ), .B(\R_DATA_TEMPR125[10] ), 
        .C(\R_DATA_TEMPR126[10] ), .D(\R_DATA_TEMPR127[10] ), .Y(
        OR4_664_Y));
    OR4 OR4_1326 (.A(\R_DATA_TEMPR96[7] ), .B(\R_DATA_TEMPR97[7] ), .C(
        \R_DATA_TEMPR98[7] ), .D(\R_DATA_TEMPR99[7] ), .Y(OR4_1326_Y));
    OR4 OR4_1348 (.A(\R_DATA_TEMPR0[35] ), .B(\R_DATA_TEMPR1[35] ), .C(
        \R_DATA_TEMPR2[35] ), .D(\R_DATA_TEMPR3[35] ), .Y(OR4_1348_Y));
    CFG3 #( .INIT(8'h4) )  CFG3_14 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_14_Y));
    OR4 OR4_623 (.A(\R_DATA_TEMPR80[17] ), .B(\R_DATA_TEMPR81[17] ), 
        .C(\R_DATA_TEMPR82[17] ), .D(\R_DATA_TEMPR83[17] ), .Y(
        OR4_623_Y));
    OR4 OR4_1621 (.A(\R_DATA_TEMPR12[17] ), .B(\R_DATA_TEMPR13[17] ), 
        .C(\R_DATA_TEMPR14[17] ), .D(\R_DATA_TEMPR15[17] ), .Y(
        OR4_1621_Y));
    OR4 OR4_1409 (.A(\R_DATA_TEMPR92[27] ), .B(\R_DATA_TEMPR93[27] ), 
        .C(\R_DATA_TEMPR94[27] ), .D(\R_DATA_TEMPR95[27] ), .Y(
        OR4_1409_Y));
    OR4 OR4_1389 (.A(\R_DATA_TEMPR80[7] ), .B(\R_DATA_TEMPR81[7] ), .C(
        \R_DATA_TEMPR82[7] ), .D(\R_DATA_TEMPR83[7] ), .Y(OR4_1389_Y));
    OR4 OR4_586 (.A(\R_DATA_TEMPR112[25] ), .B(\R_DATA_TEMPR113[25] ), 
        .C(\R_DATA_TEMPR114[25] ), .D(\R_DATA_TEMPR115[25] ), .Y(
        OR4_586_Y));
    OR4 OR4_1620 (.A(\R_DATA_TEMPR40[7] ), .B(\R_DATA_TEMPR41[7] ), .C(
        \R_DATA_TEMPR42[7] ), .D(\R_DATA_TEMPR43[7] ), .Y(OR4_1620_Y));
    OR4 OR4_1080 (.A(\R_DATA_TEMPR40[36] ), .B(\R_DATA_TEMPR41[36] ), 
        .C(\R_DATA_TEMPR42[36] ), .D(\R_DATA_TEMPR43[36] ), .Y(
        OR4_1080_Y));
    OR4 OR4_1134 (.A(\R_DATA_TEMPR108[39] ), .B(\R_DATA_TEMPR109[39] ), 
        .C(\R_DATA_TEMPR110[39] ), .D(\R_DATA_TEMPR111[39] ), .Y(
        OR4_1134_Y));
    OR4 OR4_200 (.A(\R_DATA_TEMPR120[4] ), .B(\R_DATA_TEMPR121[4] ), 
        .C(\R_DATA_TEMPR122[4] ), .D(\R_DATA_TEMPR123[4] ), .Y(
        OR4_200_Y));
    OR4 OR4_1064 (.A(OR4_102_Y), .B(OR4_1115_Y), .C(OR4_1378_Y), .D(
        OR4_328_Y), .Y(OR4_1064_Y));
    OR4 OR4_507 (.A(\R_DATA_TEMPR12[16] ), .B(\R_DATA_TEMPR13[16] ), 
        .C(\R_DATA_TEMPR14[16] ), .D(\R_DATA_TEMPR15[16] ), .Y(
        OR4_507_Y));
    OR4 OR4_1530 (.A(\R_DATA_TEMPR60[32] ), .B(\R_DATA_TEMPR61[32] ), 
        .C(\R_DATA_TEMPR62[32] ), .D(\R_DATA_TEMPR63[32] ), .Y(
        OR4_1530_Y));
    OR4 OR4_1049 (.A(\R_DATA_TEMPR12[13] ), .B(\R_DATA_TEMPR13[13] ), 
        .C(\R_DATA_TEMPR14[13] ), .D(\R_DATA_TEMPR15[13] ), .Y(
        OR4_1049_Y));
    OR4 OR4_270 (.A(\R_DATA_TEMPR88[10] ), .B(\R_DATA_TEMPR89[10] ), 
        .C(\R_DATA_TEMPR90[10] ), .D(\R_DATA_TEMPR91[10] ), .Y(
        OR4_270_Y));
    OR4 OR4_1363 (.A(\R_DATA_TEMPR4[16] ), .B(\R_DATA_TEMPR5[16] ), .C(
        \R_DATA_TEMPR6[16] ), .D(\R_DATA_TEMPR7[16] ), .Y(OR4_1363_Y));
    OR4 OR4_1170 (.A(\R_DATA_TEMPR36[18] ), .B(\R_DATA_TEMPR37[18] ), 
        .C(\R_DATA_TEMPR38[18] ), .D(\R_DATA_TEMPR39[18] ), .Y(
        OR4_1170_Y));
    OR4 OR4_929 (.A(OR4_699_Y), .B(OR4_385_Y), .C(OR4_801_Y), .D(
        OR4_629_Y), .Y(OR4_929_Y));
    OR4 OR4_920 (.A(\R_DATA_TEMPR60[36] ), .B(\R_DATA_TEMPR61[36] ), 
        .C(\R_DATA_TEMPR62[36] ), .D(\R_DATA_TEMPR63[36] ), .Y(
        OR4_920_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%106%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R106C0 (.A_DOUT({
        \R_DATA_TEMPR106[39] , \R_DATA_TEMPR106[38] , 
        \R_DATA_TEMPR106[37] , \R_DATA_TEMPR106[36] , 
        \R_DATA_TEMPR106[35] , \R_DATA_TEMPR106[34] , 
        \R_DATA_TEMPR106[33] , \R_DATA_TEMPR106[32] , 
        \R_DATA_TEMPR106[31] , \R_DATA_TEMPR106[30] , 
        \R_DATA_TEMPR106[29] , \R_DATA_TEMPR106[28] , 
        \R_DATA_TEMPR106[27] , \R_DATA_TEMPR106[26] , 
        \R_DATA_TEMPR106[25] , \R_DATA_TEMPR106[24] , 
        \R_DATA_TEMPR106[23] , \R_DATA_TEMPR106[22] , 
        \R_DATA_TEMPR106[21] , \R_DATA_TEMPR106[20] }), .B_DOUT({
        \R_DATA_TEMPR106[19] , \R_DATA_TEMPR106[18] , 
        \R_DATA_TEMPR106[17] , \R_DATA_TEMPR106[16] , 
        \R_DATA_TEMPR106[15] , \R_DATA_TEMPR106[14] , 
        \R_DATA_TEMPR106[13] , \R_DATA_TEMPR106[12] , 
        \R_DATA_TEMPR106[11] , \R_DATA_TEMPR106[10] , 
        \R_DATA_TEMPR106[9] , \R_DATA_TEMPR106[8] , 
        \R_DATA_TEMPR106[7] , \R_DATA_TEMPR106[6] , 
        \R_DATA_TEMPR106[5] , \R_DATA_TEMPR106[4] , 
        \R_DATA_TEMPR106[3] , \R_DATA_TEMPR106[2] , 
        \R_DATA_TEMPR106[1] , \R_DATA_TEMPR106[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[106][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[26] , R_ADDR[10], \BLKY0[0] }), 
        .A_CLK(CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], 
        W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], 
        W_DATA[31], W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], 
        W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], 
        W_DATA[21], W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], 
        WBYTE_EN[2]}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], 
        W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], 
        W_ADDR[0], GND, GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[26] , 
        W_ADDR[10], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA[19], 
        W_DATA[18], W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], 
        W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], W_DATA[9], 
        W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], 
        W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_890 (.A(OR4_249_Y), .B(OR4_72_Y), .C(OR4_1100_Y), .D(
        OR4_1630_Y), .Y(OR4_890_Y));
    OR4 OR4_577 (.A(OR4_284_Y), .B(OR4_1594_Y), .C(OR4_1562_Y), .D(
        OR4_705_Y), .Y(OR4_577_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[12]  (.A(CFG3_18_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[12] ));
    OR4 OR4_957 (.A(\R_DATA_TEMPR88[3] ), .B(\R_DATA_TEMPR89[3] ), .C(
        \R_DATA_TEMPR90[3] ), .D(\R_DATA_TEMPR91[3] ), .Y(OR4_957_Y));
    OR4 OR4_739 (.A(\R_DATA_TEMPR92[0] ), .B(\R_DATA_TEMPR93[0] ), .C(
        \R_DATA_TEMPR94[0] ), .D(\R_DATA_TEMPR95[0] ), .Y(OR4_739_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[21]  (.A(CFG3_22_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[21] ));
    OR4 OR4_541 (.A(\R_DATA_TEMPR52[19] ), .B(\R_DATA_TEMPR53[19] ), 
        .C(\R_DATA_TEMPR54[19] ), .D(\R_DATA_TEMPR55[19] ), .Y(
        OR4_541_Y));
    OR4 OR4_192 (.A(OR4_891_Y), .B(OR4_1345_Y), .C(OR4_671_Y), .D(
        OR4_978_Y), .Y(OR4_192_Y));
    OR4 OR4_319 (.A(OR4_779_Y), .B(OR4_798_Y), .C(OR4_780_Y), .D(
        OR4_468_Y), .Y(OR4_319_Y));
    OR4 OR4_1489 (.A(\R_DATA_TEMPR12[2] ), .B(\R_DATA_TEMPR13[2] ), .C(
        \R_DATA_TEMPR14[2] ), .D(\R_DATA_TEMPR15[2] ), .Y(OR4_1489_Y));
    OR4 OR4_1238 (.A(\R_DATA_TEMPR120[38] ), .B(\R_DATA_TEMPR121[38] ), 
        .C(\R_DATA_TEMPR122[38] ), .D(\R_DATA_TEMPR123[38] ), .Y(
        OR4_1238_Y));
    OR4 OR4_609 (.A(\R_DATA_TEMPR20[10] ), .B(\R_DATA_TEMPR21[10] ), 
        .C(\R_DATA_TEMPR22[10] ), .D(\R_DATA_TEMPR23[10] ), .Y(
        OR4_609_Y));
    OR4 OR4_1428 (.A(OR4_1142_Y), .B(OR4_1503_Y), .C(OR4_42_Y), .D(
        OR4_1236_Y), .Y(OR4_1428_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%79%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R79C0 (.A_DOUT({
        \R_DATA_TEMPR79[39] , \R_DATA_TEMPR79[38] , 
        \R_DATA_TEMPR79[37] , \R_DATA_TEMPR79[36] , 
        \R_DATA_TEMPR79[35] , \R_DATA_TEMPR79[34] , 
        \R_DATA_TEMPR79[33] , \R_DATA_TEMPR79[32] , 
        \R_DATA_TEMPR79[31] , \R_DATA_TEMPR79[30] , 
        \R_DATA_TEMPR79[29] , \R_DATA_TEMPR79[28] , 
        \R_DATA_TEMPR79[27] , \R_DATA_TEMPR79[26] , 
        \R_DATA_TEMPR79[25] , \R_DATA_TEMPR79[24] , 
        \R_DATA_TEMPR79[23] , \R_DATA_TEMPR79[22] , 
        \R_DATA_TEMPR79[21] , \R_DATA_TEMPR79[20] }), .B_DOUT({
        \R_DATA_TEMPR79[19] , \R_DATA_TEMPR79[18] , 
        \R_DATA_TEMPR79[17] , \R_DATA_TEMPR79[16] , 
        \R_DATA_TEMPR79[15] , \R_DATA_TEMPR79[14] , 
        \R_DATA_TEMPR79[13] , \R_DATA_TEMPR79[12] , 
        \R_DATA_TEMPR79[11] , \R_DATA_TEMPR79[10] , 
        \R_DATA_TEMPR79[9] , \R_DATA_TEMPR79[8] , \R_DATA_TEMPR79[7] , 
        \R_DATA_TEMPR79[6] , \R_DATA_TEMPR79[5] , \R_DATA_TEMPR79[4] , 
        \R_DATA_TEMPR79[3] , \R_DATA_TEMPR79[2] , \R_DATA_TEMPR79[1] , 
        \R_DATA_TEMPR79[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[79][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[19] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[19] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_995 (.A(\R_DATA_TEMPR44[21] ), .B(\R_DATA_TEMPR45[21] ), 
        .C(\R_DATA_TEMPR46[21] ), .D(\R_DATA_TEMPR47[21] ), .Y(
        OR4_995_Y));
    OR4 OR4_123 (.A(OR4_658_Y), .B(OR4_913_Y), .C(OR4_1104_Y), .D(
        OR4_746_Y), .Y(OR4_123_Y));
    OR4 OR4_834 (.A(\R_DATA_TEMPR68[26] ), .B(\R_DATA_TEMPR69[26] ), 
        .C(\R_DATA_TEMPR70[26] ), .D(\R_DATA_TEMPR71[26] ), .Y(
        OR4_834_Y));
    OR4 OR4_679 (.A(OR4_712_Y), .B(OR4_460_Y), .C(OR4_162_Y), .D(
        OR4_822_Y), .Y(OR4_679_Y));
    OR4 OR4_1257 (.A(\R_DATA_TEMPR24[37] ), .B(\R_DATA_TEMPR25[37] ), 
        .C(\R_DATA_TEMPR26[37] ), .D(\R_DATA_TEMPR27[37] ), .Y(
        OR4_1257_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[2]  (.A(CFG3_14_Y), .B(
        CFG3_12_Y), .Y(\BLKX2[2] ));
    OR4 OR4_206 (.A(\R_DATA_TEMPR28[33] ), .B(\R_DATA_TEMPR29[33] ), 
        .C(\R_DATA_TEMPR30[33] ), .D(\R_DATA_TEMPR31[33] ), .Y(
        OR4_206_Y));
    OR4 OR4_533 (.A(OR4_765_Y), .B(OR4_1068_Y), .C(OR4_1328_Y), .D(
        OR4_1116_Y), .Y(OR4_533_Y));
    OR4 OR4_70 (.A(\R_DATA_TEMPR40[2] ), .B(\R_DATA_TEMPR41[2] ), .C(
        \R_DATA_TEMPR42[2] ), .D(\R_DATA_TEMPR43[2] ), .Y(OR4_70_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%89%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R89C0 (.A_DOUT({
        \R_DATA_TEMPR89[39] , \R_DATA_TEMPR89[38] , 
        \R_DATA_TEMPR89[37] , \R_DATA_TEMPR89[36] , 
        \R_DATA_TEMPR89[35] , \R_DATA_TEMPR89[34] , 
        \R_DATA_TEMPR89[33] , \R_DATA_TEMPR89[32] , 
        \R_DATA_TEMPR89[31] , \R_DATA_TEMPR89[30] , 
        \R_DATA_TEMPR89[29] , \R_DATA_TEMPR89[28] , 
        \R_DATA_TEMPR89[27] , \R_DATA_TEMPR89[26] , 
        \R_DATA_TEMPR89[25] , \R_DATA_TEMPR89[24] , 
        \R_DATA_TEMPR89[23] , \R_DATA_TEMPR89[22] , 
        \R_DATA_TEMPR89[21] , \R_DATA_TEMPR89[20] }), .B_DOUT({
        \R_DATA_TEMPR89[19] , \R_DATA_TEMPR89[18] , 
        \R_DATA_TEMPR89[17] , \R_DATA_TEMPR89[16] , 
        \R_DATA_TEMPR89[15] , \R_DATA_TEMPR89[14] , 
        \R_DATA_TEMPR89[13] , \R_DATA_TEMPR89[12] , 
        \R_DATA_TEMPR89[11] , \R_DATA_TEMPR89[10] , 
        \R_DATA_TEMPR89[9] , \R_DATA_TEMPR89[8] , \R_DATA_TEMPR89[7] , 
        \R_DATA_TEMPR89[6] , \R_DATA_TEMPR89[5] , \R_DATA_TEMPR89[4] , 
        \R_DATA_TEMPR89[3] , \R_DATA_TEMPR89[2] , \R_DATA_TEMPR89[1] , 
        \R_DATA_TEMPR89[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[89][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[22] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[22] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_588 (.A(\R_DATA_TEMPR60[19] ), .B(\R_DATA_TEMPR61[19] ), 
        .C(\R_DATA_TEMPR62[19] ), .D(\R_DATA_TEMPR63[19] ), .Y(
        OR4_588_Y));
    OR4 OR4_58 (.A(\R_DATA_TEMPR12[34] ), .B(\R_DATA_TEMPR13[34] ), .C(
        \R_DATA_TEMPR14[34] ), .D(\R_DATA_TEMPR15[34] ), .Y(OR4_58_Y));
    OR4 OR4_1112 (.A(\R_DATA_TEMPR88[37] ), .B(\R_DATA_TEMPR89[37] ), 
        .C(\R_DATA_TEMPR90[37] ), .D(\R_DATA_TEMPR91[37] ), .Y(
        OR4_1112_Y));
    OR4 OR4_276 (.A(\R_DATA_TEMPR72[38] ), .B(\R_DATA_TEMPR73[38] ), 
        .C(\R_DATA_TEMPR74[38] ), .D(\R_DATA_TEMPR75[38] ), .Y(
        OR4_276_Y));
    OR4 OR4_1400 (.A(\R_DATA_TEMPR36[38] ), .B(\R_DATA_TEMPR37[38] ), 
        .C(\R_DATA_TEMPR38[38] ), .D(\R_DATA_TEMPR39[38] ), .Y(
        OR4_1400_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%63%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R63C0 (.A_DOUT({
        \R_DATA_TEMPR63[39] , \R_DATA_TEMPR63[38] , 
        \R_DATA_TEMPR63[37] , \R_DATA_TEMPR63[36] , 
        \R_DATA_TEMPR63[35] , \R_DATA_TEMPR63[34] , 
        \R_DATA_TEMPR63[33] , \R_DATA_TEMPR63[32] , 
        \R_DATA_TEMPR63[31] , \R_DATA_TEMPR63[30] , 
        \R_DATA_TEMPR63[29] , \R_DATA_TEMPR63[28] , 
        \R_DATA_TEMPR63[27] , \R_DATA_TEMPR63[26] , 
        \R_DATA_TEMPR63[25] , \R_DATA_TEMPR63[24] , 
        \R_DATA_TEMPR63[23] , \R_DATA_TEMPR63[22] , 
        \R_DATA_TEMPR63[21] , \R_DATA_TEMPR63[20] }), .B_DOUT({
        \R_DATA_TEMPR63[19] , \R_DATA_TEMPR63[18] , 
        \R_DATA_TEMPR63[17] , \R_DATA_TEMPR63[16] , 
        \R_DATA_TEMPR63[15] , \R_DATA_TEMPR63[14] , 
        \R_DATA_TEMPR63[13] , \R_DATA_TEMPR63[12] , 
        \R_DATA_TEMPR63[11] , \R_DATA_TEMPR63[10] , 
        \R_DATA_TEMPR63[9] , \R_DATA_TEMPR63[8] , \R_DATA_TEMPR63[7] , 
        \R_DATA_TEMPR63[6] , \R_DATA_TEMPR63[5] , \R_DATA_TEMPR63[4] , 
        \R_DATA_TEMPR63[3] , \R_DATA_TEMPR63[2] , \R_DATA_TEMPR63[1] , 
        \R_DATA_TEMPR63[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[63][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[15] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[15] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_242 (.A(OR4_1608_Y), .B(OR4_824_Y), .C(OR4_1631_Y), .D(
        OR4_254_Y), .Y(OR4_242_Y));
    OR4 OR4_77 (.A(OR4_332_Y), .B(OR4_308_Y), .C(OR4_270_Y), .D(
        OR4_1041_Y), .Y(OR4_77_Y));
    OR4 OR4_1456 (.A(OR4_482_Y), .B(OR4_788_Y), .C(OR4_1021_Y), .D(
        OR4_839_Y), .Y(OR4_1456_Y));
    OR4 OR4_1370 (.A(\R_DATA_TEMPR24[25] ), .B(\R_DATA_TEMPR25[25] ), 
        .C(\R_DATA_TEMPR26[25] ), .D(\R_DATA_TEMPR27[25] ), .Y(
        OR4_1370_Y));
    OR4 OR4_1354 (.A(OR4_1292_Y), .B(OR4_1280_Y), .C(OR4_1169_Y), .D(
        OR4_1582_Y), .Y(OR4_1354_Y));
    OR4 OR4_604 (.A(\R_DATA_TEMPR44[34] ), .B(\R_DATA_TEMPR45[34] ), 
        .C(\R_DATA_TEMPR46[34] ), .D(\R_DATA_TEMPR47[34] ), .Y(
        OR4_604_Y));
    OR4 OR4_1124 (.A(OR4_905_Y), .B(OR4_931_Y), .C(OR4_909_Y), .D(
        OR4_62_Y), .Y(OR4_1124_Y));
    OR4 OR4_299 (.A(\R_DATA_TEMPR24[39] ), .B(\R_DATA_TEMPR25[39] ), 
        .C(\R_DATA_TEMPR26[39] ), .D(\R_DATA_TEMPR27[39] ), .Y(
        OR4_299_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[16]  (.A(CFG3_13_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[16] ));
    OR4 OR4_1094 (.A(\R_DATA_TEMPR28[25] ), .B(\R_DATA_TEMPR29[25] ), 
        .C(\R_DATA_TEMPR30[25] ), .D(\R_DATA_TEMPR31[25] ), .Y(
        OR4_1094_Y));
    OR4 OR4_1101 (.A(\R_DATA_TEMPR16[20] ), .B(\R_DATA_TEMPR17[20] ), 
        .C(\R_DATA_TEMPR18[20] ), .D(\R_DATA_TEMPR19[20] ), .Y(
        OR4_1101_Y));
    OR4 OR4_674 (.A(\R_DATA_TEMPR56[11] ), .B(\R_DATA_TEMPR57[11] ), 
        .C(\R_DATA_TEMPR58[11] ), .D(\R_DATA_TEMPR59[11] ), .Y(
        OR4_674_Y));
    OR4 OR4_455 (.A(OR4_1495_Y), .B(OR4_147_Y), .C(OR4_1244_Y), .D(
        OR4_469_Y), .Y(OR4_455_Y));
    OR4 OR4_1520 (.A(\R_DATA_TEMPR52[30] ), .B(\R_DATA_TEMPR53[30] ), 
        .C(\R_DATA_TEMPR54[30] ), .D(\R_DATA_TEMPR55[30] ), .Y(
        OR4_1520_Y));
    OR4 OR4_486 (.A(OR4_65_Y), .B(OR4_845_Y), .C(OR4_1316_Y), .D(
        OR4_1621_Y), .Y(OR4_486_Y));
    OR4 OR4_1393 (.A(OR4_228_Y), .B(OR4_30_Y), .C(OR4_1308_Y), .D(
        OR4_1127_Y), .Y(OR4_1393_Y));
    OR4 \OR4_R_DATA[5]  (.A(OR4_269_Y), .B(OR4_1553_Y), .C(OR4_1029_Y), 
        .D(OR4_1358_Y), .Y(R_DATA[5]));
    OR4 OR4_340 (.A(\R_DATA_TEMPR76[6] ), .B(\R_DATA_TEMPR77[6] ), .C(
        \R_DATA_TEMPR78[6] ), .D(\R_DATA_TEMPR79[6] ), .Y(OR4_340_Y));
    OR4 OR4_1066 (.A(\R_DATA_TEMPR64[12] ), .B(\R_DATA_TEMPR65[12] ), 
        .C(\R_DATA_TEMPR66[12] ), .D(\R_DATA_TEMPR67[12] ), .Y(
        OR4_1066_Y));
    OR4 OR4_1506 (.A(\R_DATA_TEMPR4[19] ), .B(\R_DATA_TEMPR5[19] ), .C(
        \R_DATA_TEMPR6[19] ), .D(\R_DATA_TEMPR7[19] ), .Y(OR4_1506_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%75%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R75C0 (.A_DOUT({
        \R_DATA_TEMPR75[39] , \R_DATA_TEMPR75[38] , 
        \R_DATA_TEMPR75[37] , \R_DATA_TEMPR75[36] , 
        \R_DATA_TEMPR75[35] , \R_DATA_TEMPR75[34] , 
        \R_DATA_TEMPR75[33] , \R_DATA_TEMPR75[32] , 
        \R_DATA_TEMPR75[31] , \R_DATA_TEMPR75[30] , 
        \R_DATA_TEMPR75[29] , \R_DATA_TEMPR75[28] , 
        \R_DATA_TEMPR75[27] , \R_DATA_TEMPR75[26] , 
        \R_DATA_TEMPR75[25] , \R_DATA_TEMPR75[24] , 
        \R_DATA_TEMPR75[23] , \R_DATA_TEMPR75[22] , 
        \R_DATA_TEMPR75[21] , \R_DATA_TEMPR75[20] }), .B_DOUT({
        \R_DATA_TEMPR75[19] , \R_DATA_TEMPR75[18] , 
        \R_DATA_TEMPR75[17] , \R_DATA_TEMPR75[16] , 
        \R_DATA_TEMPR75[15] , \R_DATA_TEMPR75[14] , 
        \R_DATA_TEMPR75[13] , \R_DATA_TEMPR75[12] , 
        \R_DATA_TEMPR75[11] , \R_DATA_TEMPR75[10] , 
        \R_DATA_TEMPR75[9] , \R_DATA_TEMPR75[8] , \R_DATA_TEMPR75[7] , 
        \R_DATA_TEMPR75[6] , \R_DATA_TEMPR75[5] , \R_DATA_TEMPR75[4] , 
        \R_DATA_TEMPR75[3] , \R_DATA_TEMPR75[2] , \R_DATA_TEMPR75[1] , 
        \R_DATA_TEMPR75[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[75][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[18] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[18] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1639 (.A(\R_DATA_TEMPR92[32] ), .B(\R_DATA_TEMPR93[32] ), 
        .C(\R_DATA_TEMPR94[32] ), .D(\R_DATA_TEMPR95[32] ), .Y(
        OR4_1639_Y));
    OR4 OR4_1135 (.A(\R_DATA_TEMPR24[8] ), .B(\R_DATA_TEMPR25[8] ), .C(
        \R_DATA_TEMPR26[8] ), .D(\R_DATA_TEMPR27[8] ), .Y(OR4_1135_Y));
    OR4 OR4_719 (.A(\R_DATA_TEMPR72[18] ), .B(\R_DATA_TEMPR73[18] ), 
        .C(\R_DATA_TEMPR74[18] ), .D(\R_DATA_TEMPR75[18] ), .Y(
        OR4_719_Y));
    OR4 OR4_1228 (.A(\R_DATA_TEMPR80[33] ), .B(\R_DATA_TEMPR81[33] ), 
        .C(\R_DATA_TEMPR82[33] ), .D(\R_DATA_TEMPR83[33] ), .Y(
        OR4_1228_Y));
    OR4 OR4_820 (.A(OR4_216_Y), .B(OR2_30_Y), .C(\R_DATA_TEMPR86[20] ), 
        .D(\R_DATA_TEMPR87[20] ), .Y(OR4_820_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%54%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R54C0 (.A_DOUT({
        \R_DATA_TEMPR54[39] , \R_DATA_TEMPR54[38] , 
        \R_DATA_TEMPR54[37] , \R_DATA_TEMPR54[36] , 
        \R_DATA_TEMPR54[35] , \R_DATA_TEMPR54[34] , 
        \R_DATA_TEMPR54[33] , \R_DATA_TEMPR54[32] , 
        \R_DATA_TEMPR54[31] , \R_DATA_TEMPR54[30] , 
        \R_DATA_TEMPR54[29] , \R_DATA_TEMPR54[28] , 
        \R_DATA_TEMPR54[27] , \R_DATA_TEMPR54[26] , 
        \R_DATA_TEMPR54[25] , \R_DATA_TEMPR54[24] , 
        \R_DATA_TEMPR54[23] , \R_DATA_TEMPR54[22] , 
        \R_DATA_TEMPR54[21] , \R_DATA_TEMPR54[20] }), .B_DOUT({
        \R_DATA_TEMPR54[19] , \R_DATA_TEMPR54[18] , 
        \R_DATA_TEMPR54[17] , \R_DATA_TEMPR54[16] , 
        \R_DATA_TEMPR54[15] , \R_DATA_TEMPR54[14] , 
        \R_DATA_TEMPR54[13] , \R_DATA_TEMPR54[12] , 
        \R_DATA_TEMPR54[11] , \R_DATA_TEMPR54[10] , 
        \R_DATA_TEMPR54[9] , \R_DATA_TEMPR54[8] , \R_DATA_TEMPR54[7] , 
        \R_DATA_TEMPR54[6] , \R_DATA_TEMPR54[5] , \R_DATA_TEMPR54[4] , 
        \R_DATA_TEMPR54[3] , \R_DATA_TEMPR54[2] , \R_DATA_TEMPR54[1] , 
        \R_DATA_TEMPR54[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[54][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[13] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[13] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1480 (.A(\R_DATA_TEMPR24[38] ), .B(\R_DATA_TEMPR25[38] ), 
        .C(\R_DATA_TEMPR26[38] ), .D(\R_DATA_TEMPR27[38] ), .Y(
        OR4_1480_Y));
    OR4 OR4_1031 (.A(\R_DATA_TEMPR16[26] ), .B(\R_DATA_TEMPR17[26] ), 
        .C(\R_DATA_TEMPR18[26] ), .D(\R_DATA_TEMPR19[26] ), .Y(
        OR4_1031_Y));
    OR4 OR4_899 (.A(OR4_1550_Y), .B(OR4_467_Y), .C(OR4_1156_Y), .D(
        OR4_202_Y), .Y(OR4_899_Y));
    OR4 \OR4_R_DATA[11]  (.A(OR4_2_Y), .B(OR4_1560_Y), .C(OR4_1590_Y), 
        .D(OR4_1078_Y), .Y(R_DATA[11]));
    OR4 OR4_122 (.A(\R_DATA_TEMPR40[15] ), .B(\R_DATA_TEMPR41[15] ), 
        .C(\R_DATA_TEMPR42[15] ), .D(\R_DATA_TEMPR43[15] ), .Y(
        OR4_122_Y));
    OR4 OR4_1361 (.A(\R_DATA_TEMPR96[12] ), .B(\R_DATA_TEMPR97[12] ), 
        .C(\R_DATA_TEMPR98[12] ), .D(\R_DATA_TEMPR99[12] ), .Y(
        OR4_1361_Y));
    OR4 OR4_843 (.A(OR4_535_Y), .B(OR4_781_Y), .C(OR4_967_Y), .D(
        OR4_884_Y), .Y(OR4_843_Y));
    OR4 OR4_814 (.A(OR4_1022_Y), .B(OR4_542_Y), .C(OR4_595_Y), .D(
        OR4_966_Y), .Y(OR4_814_Y));
    OR4 OR4_382 (.A(\R_DATA_TEMPR104[5] ), .B(\R_DATA_TEMPR105[5] ), 
        .C(\R_DATA_TEMPR106[5] ), .D(\R_DATA_TEMPR107[5] ), .Y(
        OR4_382_Y));
    OR4 OR4_925 (.A(OR4_1406_Y), .B(OR4_1214_Y), .C(OR4_614_Y), .D(
        OR4_1126_Y), .Y(OR4_925_Y));
    OR4 \OR4_R_DATA[9]  (.A(OR4_219_Y), .B(OR4_529_Y), .C(OR4_939_Y), 
        .D(OR4_1259_Y), .Y(R_DATA[9]));
    OR4 OR4_1359 (.A(OR4_947_Y), .B(OR2_0_Y), .C(\R_DATA_TEMPR86[16] ), 
        .D(\R_DATA_TEMPR87[16] ), .Y(OR4_1359_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%44%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R44C0 (.A_DOUT({
        \R_DATA_TEMPR44[39] , \R_DATA_TEMPR44[38] , 
        \R_DATA_TEMPR44[37] , \R_DATA_TEMPR44[36] , 
        \R_DATA_TEMPR44[35] , \R_DATA_TEMPR44[34] , 
        \R_DATA_TEMPR44[33] , \R_DATA_TEMPR44[32] , 
        \R_DATA_TEMPR44[31] , \R_DATA_TEMPR44[30] , 
        \R_DATA_TEMPR44[29] , \R_DATA_TEMPR44[28] , 
        \R_DATA_TEMPR44[27] , \R_DATA_TEMPR44[26] , 
        \R_DATA_TEMPR44[25] , \R_DATA_TEMPR44[24] , 
        \R_DATA_TEMPR44[23] , \R_DATA_TEMPR44[22] , 
        \R_DATA_TEMPR44[21] , \R_DATA_TEMPR44[20] }), .B_DOUT({
        \R_DATA_TEMPR44[19] , \R_DATA_TEMPR44[18] , 
        \R_DATA_TEMPR44[17] , \R_DATA_TEMPR44[16] , 
        \R_DATA_TEMPR44[15] , \R_DATA_TEMPR44[14] , 
        \R_DATA_TEMPR44[13] , \R_DATA_TEMPR44[12] , 
        \R_DATA_TEMPR44[11] , \R_DATA_TEMPR44[10] , 
        \R_DATA_TEMPR44[9] , \R_DATA_TEMPR44[8] , \R_DATA_TEMPR44[7] , 
        \R_DATA_TEMPR44[6] , \R_DATA_TEMPR44[5] , \R_DATA_TEMPR44[4] , 
        \R_DATA_TEMPR44[3] , \R_DATA_TEMPR44[2] , \R_DATA_TEMPR44[1] , 
        \R_DATA_TEMPR44[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[44][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[11] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[11] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%85%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R85C0 (.A_DOUT({
        \R_DATA_TEMPR85[39] , \R_DATA_TEMPR85[38] , 
        \R_DATA_TEMPR85[37] , \R_DATA_TEMPR85[36] , 
        \R_DATA_TEMPR85[35] , \R_DATA_TEMPR85[34] , 
        \R_DATA_TEMPR85[33] , \R_DATA_TEMPR85[32] , 
        \R_DATA_TEMPR85[31] , \R_DATA_TEMPR85[30] , 
        \R_DATA_TEMPR85[29] , \R_DATA_TEMPR85[28] , 
        \R_DATA_TEMPR85[27] , \R_DATA_TEMPR85[26] , 
        \R_DATA_TEMPR85[25] , \R_DATA_TEMPR85[24] , 
        \R_DATA_TEMPR85[23] , \R_DATA_TEMPR85[22] , 
        \R_DATA_TEMPR85[21] , \R_DATA_TEMPR85[20] }), .B_DOUT({
        \R_DATA_TEMPR85[19] , \R_DATA_TEMPR85[18] , 
        \R_DATA_TEMPR85[17] , \R_DATA_TEMPR85[16] , 
        \R_DATA_TEMPR85[15] , \R_DATA_TEMPR85[14] , 
        \R_DATA_TEMPR85[13] , \R_DATA_TEMPR85[12] , 
        \R_DATA_TEMPR85[11] , \R_DATA_TEMPR85[10] , 
        \R_DATA_TEMPR85[9] , \R_DATA_TEMPR85[8] , \R_DATA_TEMPR85[7] , 
        \R_DATA_TEMPR85[6] , \R_DATA_TEMPR85[5] , \R_DATA_TEMPR85[4] , 
        \R_DATA_TEMPR85[3] , \R_DATA_TEMPR85[2] , \R_DATA_TEMPR85[1] , 
        \R_DATA_TEMPR85[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[85][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[21] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[21] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_18 (.A(\R_DATA_TEMPR44[35] ), .B(\R_DATA_TEMPR45[35] ), .C(
        \R_DATA_TEMPR46[35] ), .D(\R_DATA_TEMPR47[35] ), .Y(OR4_18_Y));
    OR4 OR4_513 (.A(\R_DATA_TEMPR104[3] ), .B(\R_DATA_TEMPR105[3] ), 
        .C(\R_DATA_TEMPR106[3] ), .D(\R_DATA_TEMPR107[3] ), .Y(
        OR4_513_Y));
    OR4 OR4_34 (.A(\R_DATA_TEMPR20[12] ), .B(\R_DATA_TEMPR21[12] ), .C(
        \R_DATA_TEMPR22[12] ), .D(\R_DATA_TEMPR23[12] ), .Y(OR4_34_Y));
    OR4 OR4_1181 (.A(\R_DATA_TEMPR28[31] ), .B(\R_DATA_TEMPR29[31] ), 
        .C(\R_DATA_TEMPR30[31] ), .D(\R_DATA_TEMPR31[31] ), .Y(
        OR4_1181_Y));
    OR4 OR4_1050 (.A(\R_DATA_TEMPR52[20] ), .B(\R_DATA_TEMPR53[20] ), 
        .C(\R_DATA_TEMPR54[20] ), .D(\R_DATA_TEMPR55[20] ), .Y(
        OR4_1050_Y));
    OR4 OR4_1147 (.A(\R_DATA_TEMPR0[22] ), .B(\R_DATA_TEMPR1[22] ), .C(
        \R_DATA_TEMPR2[22] ), .D(\R_DATA_TEMPR3[22] ), .Y(OR4_1147_Y));
    OR4 OR4_1407 (.A(\R_DATA_TEMPR32[2] ), .B(\R_DATA_TEMPR33[2] ), .C(
        \R_DATA_TEMPR34[2] ), .D(\R_DATA_TEMPR35[2] ), .Y(OR4_1407_Y));
    OR4 OR4_1275 (.A(\R_DATA_TEMPR76[2] ), .B(\R_DATA_TEMPR77[2] ), .C(
        \R_DATA_TEMPR78[2] ), .D(\R_DATA_TEMPR79[2] ), .Y(OR4_1275_Y));
    OR4 OR4_868 (.A(\R_DATA_TEMPR20[1] ), .B(\R_DATA_TEMPR21[1] ), .C(
        \R_DATA_TEMPR22[1] ), .D(\R_DATA_TEMPR23[1] ), .Y(OR4_868_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%93%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R93C0 (.A_DOUT({
        \R_DATA_TEMPR93[39] , \R_DATA_TEMPR93[38] , 
        \R_DATA_TEMPR93[37] , \R_DATA_TEMPR93[36] , 
        \R_DATA_TEMPR93[35] , \R_DATA_TEMPR93[34] , 
        \R_DATA_TEMPR93[33] , \R_DATA_TEMPR93[32] , 
        \R_DATA_TEMPR93[31] , \R_DATA_TEMPR93[30] , 
        \R_DATA_TEMPR93[29] , \R_DATA_TEMPR93[28] , 
        \R_DATA_TEMPR93[27] , \R_DATA_TEMPR93[26] , 
        \R_DATA_TEMPR93[25] , \R_DATA_TEMPR93[24] , 
        \R_DATA_TEMPR93[23] , \R_DATA_TEMPR93[22] , 
        \R_DATA_TEMPR93[21] , \R_DATA_TEMPR93[20] }), .B_DOUT({
        \R_DATA_TEMPR93[19] , \R_DATA_TEMPR93[18] , 
        \R_DATA_TEMPR93[17] , \R_DATA_TEMPR93[16] , 
        \R_DATA_TEMPR93[15] , \R_DATA_TEMPR93[14] , 
        \R_DATA_TEMPR93[13] , \R_DATA_TEMPR93[12] , 
        \R_DATA_TEMPR93[11] , \R_DATA_TEMPR93[10] , 
        \R_DATA_TEMPR93[9] , \R_DATA_TEMPR93[8] , \R_DATA_TEMPR93[7] , 
        \R_DATA_TEMPR93[6] , \R_DATA_TEMPR93[5] , \R_DATA_TEMPR93[4] , 
        \R_DATA_TEMPR93[3] , \R_DATA_TEMPR93[2] , \R_DATA_TEMPR93[1] , 
        \R_DATA_TEMPR93[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[93][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[23] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[23] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1571 (.A(\R_DATA_TEMPR92[29] ), .B(\R_DATA_TEMPR93[29] ), 
        .C(\R_DATA_TEMPR94[29] ), .D(\R_DATA_TEMPR95[29] ), .Y(
        OR4_1571_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%8%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C0 (.A_DOUT({
        \R_DATA_TEMPR8[39] , \R_DATA_TEMPR8[38] , \R_DATA_TEMPR8[37] , 
        \R_DATA_TEMPR8[36] , \R_DATA_TEMPR8[35] , \R_DATA_TEMPR8[34] , 
        \R_DATA_TEMPR8[33] , \R_DATA_TEMPR8[32] , \R_DATA_TEMPR8[31] , 
        \R_DATA_TEMPR8[30] , \R_DATA_TEMPR8[29] , \R_DATA_TEMPR8[28] , 
        \R_DATA_TEMPR8[27] , \R_DATA_TEMPR8[26] , \R_DATA_TEMPR8[25] , 
        \R_DATA_TEMPR8[24] , \R_DATA_TEMPR8[23] , \R_DATA_TEMPR8[22] , 
        \R_DATA_TEMPR8[21] , \R_DATA_TEMPR8[20] }), .B_DOUT({
        \R_DATA_TEMPR8[19] , \R_DATA_TEMPR8[18] , \R_DATA_TEMPR8[17] , 
        \R_DATA_TEMPR8[16] , \R_DATA_TEMPR8[15] , \R_DATA_TEMPR8[14] , 
        \R_DATA_TEMPR8[13] , \R_DATA_TEMPR8[12] , \R_DATA_TEMPR8[11] , 
        \R_DATA_TEMPR8[10] , \R_DATA_TEMPR8[9] , \R_DATA_TEMPR8[8] , 
        \R_DATA_TEMPR8[7] , \R_DATA_TEMPR8[6] , \R_DATA_TEMPR8[5] , 
        \R_DATA_TEMPR8[4] , \R_DATA_TEMPR8[3] , \R_DATA_TEMPR8[2] , 
        \R_DATA_TEMPR8[1] , \R_DATA_TEMPR8[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[8][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_454 (.A(OR4_689_Y), .B(OR4_508_Y), .C(OR4_485_Y), .D(
        OR4_152_Y), .Y(OR4_454_Y));
    OR4 OR4_1033 (.A(\R_DATA_TEMPR60[13] ), .B(\R_DATA_TEMPR61[13] ), 
        .C(\R_DATA_TEMPR62[13] ), .D(\R_DATA_TEMPR63[13] ), .Y(
        OR4_1033_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[11]  (.A(CFG3_19_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[11] ));
    OR4 OR4_1586 (.A(\R_DATA_TEMPR120[20] ), .B(\R_DATA_TEMPR121[20] ), 
        .C(\R_DATA_TEMPR122[20] ), .D(\R_DATA_TEMPR123[20] ), .Y(
        OR4_1586_Y));
    OR4 \OR4_R_DATA[35]  (.A(OR4_158_Y), .B(OR4_940_Y), .C(OR4_1579_Y), 
        .D(OR4_1111_Y), .Y(R_DATA[35]));
    OR4 OR4_1005 (.A(OR4_1392_Y), .B(OR4_393_Y), .C(OR4_919_Y), .D(
        OR4_336_Y), .Y(OR4_1005_Y));
    OR4 \OR4_R_DATA[10]  (.A(OR4_1342_Y), .B(OR4_77_Y), .C(OR4_813_Y), 
        .D(OR4_186_Y), .Y(R_DATA[10]));
    OR4 OR4_1432 (.A(\R_DATA_TEMPR36[26] ), .B(\R_DATA_TEMPR37[26] ), 
        .C(\R_DATA_TEMPR38[26] ), .D(\R_DATA_TEMPR39[26] ), .Y(
        OR4_1432_Y));
    OR4 OR4_229 (.A(OR4_106_Y), .B(OR4_562_Y), .C(OR4_1521_Y), .D(
        OR4_199_Y), .Y(OR4_229_Y));
    OR4 OR4_356 (.A(OR4_1117_Y), .B(OR4_361_Y), .C(OR4_1135_Y), .D(
        OR4_1414_Y), .Y(OR4_356_Y));
    OR4 OR4_797 (.A(\R_DATA_TEMPR96[34] ), .B(\R_DATA_TEMPR97[34] ), 
        .C(\R_DATA_TEMPR98[34] ), .D(\R_DATA_TEMPR99[34] ), .Y(
        OR4_797_Y));
    OR4 OR4_1459 (.A(\R_DATA_TEMPR52[25] ), .B(\R_DATA_TEMPR53[25] ), 
        .C(\R_DATA_TEMPR54[25] ), .D(\R_DATA_TEMPR55[25] ), .Y(
        OR4_1459_Y));
    OR4 OR4_794 (.A(\R_DATA_TEMPR112[21] ), .B(\R_DATA_TEMPR113[21] ), 
        .C(\R_DATA_TEMPR114[21] ), .D(\R_DATA_TEMPR115[21] ), .Y(
        OR4_794_Y));
    OR4 OR4_1096 (.A(OR4_120_Y), .B(OR4_443_Y), .C(OR4_674_Y), .D(
        OR4_493_Y), .Y(OR4_1096_Y));
    OR2 OR2_23 (.A(\R_DATA_TEMPR84[29] ), .B(\R_DATA_TEMPR85[29] ), .Y(
        OR2_23_Y));
    OR4 OR4_261 (.A(OR4_1552_Y), .B(OR4_1296_Y), .C(OR4_1000_Y), .D(
        OR4_1121_Y), .Y(OR4_261_Y));
    OR4 OR4_29 (.A(\R_DATA_TEMPR28[22] ), .B(\R_DATA_TEMPR29[22] ), .C(
        \R_DATA_TEMPR30[22] ), .D(\R_DATA_TEMPR31[22] ), .Y(OR4_29_Y));
    OR4 \OR4_R_DATA[16]  (.A(OR4_766_Y), .B(OR4_10_Y), .C(OR4_323_Y), 
        .D(OR4_395_Y), .Y(R_DATA[16]));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%108%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R108C0 (.A_DOUT({
        \R_DATA_TEMPR108[39] , \R_DATA_TEMPR108[38] , 
        \R_DATA_TEMPR108[37] , \R_DATA_TEMPR108[36] , 
        \R_DATA_TEMPR108[35] , \R_DATA_TEMPR108[34] , 
        \R_DATA_TEMPR108[33] , \R_DATA_TEMPR108[32] , 
        \R_DATA_TEMPR108[31] , \R_DATA_TEMPR108[30] , 
        \R_DATA_TEMPR108[29] , \R_DATA_TEMPR108[28] , 
        \R_DATA_TEMPR108[27] , \R_DATA_TEMPR108[26] , 
        \R_DATA_TEMPR108[25] , \R_DATA_TEMPR108[24] , 
        \R_DATA_TEMPR108[23] , \R_DATA_TEMPR108[22] , 
        \R_DATA_TEMPR108[21] , \R_DATA_TEMPR108[20] }), .B_DOUT({
        \R_DATA_TEMPR108[19] , \R_DATA_TEMPR108[18] , 
        \R_DATA_TEMPR108[17] , \R_DATA_TEMPR108[16] , 
        \R_DATA_TEMPR108[15] , \R_DATA_TEMPR108[14] , 
        \R_DATA_TEMPR108[13] , \R_DATA_TEMPR108[12] , 
        \R_DATA_TEMPR108[11] , \R_DATA_TEMPR108[10] , 
        \R_DATA_TEMPR108[9] , \R_DATA_TEMPR108[8] , 
        \R_DATA_TEMPR108[7] , \R_DATA_TEMPR108[6] , 
        \R_DATA_TEMPR108[5] , \R_DATA_TEMPR108[4] , 
        \R_DATA_TEMPR108[3] , \R_DATA_TEMPR108[2] , 
        \R_DATA_TEMPR108[1] , \R_DATA_TEMPR108[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[108][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[27] , \BLKY1[0] , \BLKY0[0] }), 
        .A_CLK(CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], 
        W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], 
        W_DATA[31], W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], 
        W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], 
        W_DATA[21], W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], 
        WBYTE_EN[2]}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], 
        W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], 
        W_ADDR[0], GND, GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[27] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA[19], 
        W_DATA[18], W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], 
        W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], W_DATA[9], 
        W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], 
        W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1629 (.A(\R_DATA_TEMPR72[7] ), .B(\R_DATA_TEMPR73[7] ), .C(
        \R_DATA_TEMPR74[7] ), .D(\R_DATA_TEMPR75[7] ), .Y(OR4_1629_Y));
    OR4 OR4_1125 (.A(\R_DATA_TEMPR92[15] ), .B(\R_DATA_TEMPR93[15] ), 
        .C(\R_DATA_TEMPR94[15] ), .D(\R_DATA_TEMPR95[15] ), .Y(
        OR4_1125_Y));
    OR4 OR4_280 (.A(\R_DATA_TEMPR64[34] ), .B(\R_DATA_TEMPR65[34] ), 
        .C(\R_DATA_TEMPR66[34] ), .D(\R_DATA_TEMPR67[34] ), .Y(
        OR4_280_Y));
    OR4 OR4_1487 (.A(\R_DATA_TEMPR120[2] ), .B(\R_DATA_TEMPR121[2] ), 
        .C(\R_DATA_TEMPR122[2] ), .D(\R_DATA_TEMPR123[2] ), .Y(
        OR4_1487_Y));
    OR4 OR4_891 (.A(\R_DATA_TEMPR0[4] ), .B(\R_DATA_TEMPR1[4] ), .C(
        \R_DATA_TEMPR2[4] ), .D(\R_DATA_TEMPR3[4] ), .Y(OR4_891_Y));
    OR4 OR4_587 (.A(OR4_730_Y), .B(OR4_985_Y), .C(OR4_505_Y), .D(
        OR4_239_Y), .Y(OR4_587_Y));
    OR4 OR4_1021 (.A(\R_DATA_TEMPR56[16] ), .B(\R_DATA_TEMPR57[16] ), 
        .C(\R_DATA_TEMPR58[16] ), .D(\R_DATA_TEMPR59[16] ), .Y(
        OR4_1021_Y));
    OR4 OR4_1391 (.A(\R_DATA_TEMPR80[18] ), .B(\R_DATA_TEMPR81[18] ), 
        .C(\R_DATA_TEMPR82[18] ), .D(\R_DATA_TEMPR83[18] ), .Y(
        OR4_1391_Y));
    OR4 OR4_545 (.A(\R_DATA_TEMPR60[37] ), .B(\R_DATA_TEMPR61[37] ), 
        .C(\R_DATA_TEMPR62[37] ), .D(\R_DATA_TEMPR63[37] ), .Y(
        OR4_545_Y));
    OR4 OR4_233 (.A(\R_DATA_TEMPR8[34] ), .B(\R_DATA_TEMPR9[34] ), .C(
        \R_DATA_TEMPR10[34] ), .D(\R_DATA_TEMPR11[34] ), .Y(OR4_233_Y));
    OR4 OR4_1085 (.A(OR4_331_Y), .B(OR4_313_Y), .C(OR4_838_Y), .D(
        OR4_234_Y), .Y(OR4_1085_Y));
    OR4 OR4_829 (.A(\R_DATA_TEMPR68[35] ), .B(\R_DATA_TEMPR69[35] ), 
        .C(\R_DATA_TEMPR70[35] ), .D(\R_DATA_TEMPR71[35] ), .Y(
        OR4_829_Y));
    OR4 OR4_562 (.A(\R_DATA_TEMPR4[6] ), .B(\R_DATA_TEMPR5[6] ), .C(
        \R_DATA_TEMPR6[6] ), .D(\R_DATA_TEMPR7[6] ), .Y(OR4_562_Y));
    OR4 OR4_689 (.A(OR4_936_Y), .B(OR4_450_Y), .C(OR4_504_Y), .D(
        OR4_981_Y), .Y(OR4_689_Y));
    OR4 OR4_643 (.A(\R_DATA_TEMPR36[8] ), .B(\R_DATA_TEMPR37[8] ), .C(
        \R_DATA_TEMPR38[8] ), .D(\R_DATA_TEMPR39[8] ), .Y(OR4_643_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%50%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R50C0 (.A_DOUT({
        \R_DATA_TEMPR50[39] , \R_DATA_TEMPR50[38] , 
        \R_DATA_TEMPR50[37] , \R_DATA_TEMPR50[36] , 
        \R_DATA_TEMPR50[35] , \R_DATA_TEMPR50[34] , 
        \R_DATA_TEMPR50[33] , \R_DATA_TEMPR50[32] , 
        \R_DATA_TEMPR50[31] , \R_DATA_TEMPR50[30] , 
        \R_DATA_TEMPR50[29] , \R_DATA_TEMPR50[28] , 
        \R_DATA_TEMPR50[27] , \R_DATA_TEMPR50[26] , 
        \R_DATA_TEMPR50[25] , \R_DATA_TEMPR50[24] , 
        \R_DATA_TEMPR50[23] , \R_DATA_TEMPR50[22] , 
        \R_DATA_TEMPR50[21] , \R_DATA_TEMPR50[20] }), .B_DOUT({
        \R_DATA_TEMPR50[19] , \R_DATA_TEMPR50[18] , 
        \R_DATA_TEMPR50[17] , \R_DATA_TEMPR50[16] , 
        \R_DATA_TEMPR50[15] , \R_DATA_TEMPR50[14] , 
        \R_DATA_TEMPR50[13] , \R_DATA_TEMPR50[12] , 
        \R_DATA_TEMPR50[11] , \R_DATA_TEMPR50[10] , 
        \R_DATA_TEMPR50[9] , \R_DATA_TEMPR50[8] , \R_DATA_TEMPR50[7] , 
        \R_DATA_TEMPR50[6] , \R_DATA_TEMPR50[5] , \R_DATA_TEMPR50[4] , 
        \R_DATA_TEMPR50[3] , \R_DATA_TEMPR50[2] , \R_DATA_TEMPR50[1] , 
        \R_DATA_TEMPR50[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[50][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[12] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[12] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_938 (.A(\R_DATA_TEMPR72[10] ), .B(\R_DATA_TEMPR73[10] ), 
        .C(\R_DATA_TEMPR74[10] ), .D(\R_DATA_TEMPR75[10] ), .Y(
        OR4_938_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[4]  (.A(CFG3_18_Y), .B(CFG3_2_Y)
        , .Y(\BLKY2[4] ));
    OR4 OR4_1240 (.A(\R_DATA_TEMPR16[32] ), .B(\R_DATA_TEMPR17[32] ), 
        .C(\R_DATA_TEMPR18[32] ), .D(\R_DATA_TEMPR19[32] ), .Y(
        OR4_1240_Y));
    OR4 OR4_1023 (.A(\R_DATA_TEMPR72[12] ), .B(\R_DATA_TEMPR73[12] ), 
        .C(\R_DATA_TEMPR74[12] ), .D(\R_DATA_TEMPR75[12] ), .Y(
        OR4_1023_Y));
    OR4 OR4_1518 (.A(\R_DATA_TEMPR40[9] ), .B(\R_DATA_TEMPR41[9] ), .C(
        \R_DATA_TEMPR42[9] ), .D(\R_DATA_TEMPR43[9] ), .Y(OR4_1518_Y));
    OR4 OR4_286 (.A(\R_DATA_TEMPR4[15] ), .B(\R_DATA_TEMPR5[15] ), .C(
        \R_DATA_TEMPR6[15] ), .D(\R_DATA_TEMPR7[15] ), .Y(OR4_286_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%40%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R40C0 (.A_DOUT({
        \R_DATA_TEMPR40[39] , \R_DATA_TEMPR40[38] , 
        \R_DATA_TEMPR40[37] , \R_DATA_TEMPR40[36] , 
        \R_DATA_TEMPR40[35] , \R_DATA_TEMPR40[34] , 
        \R_DATA_TEMPR40[33] , \R_DATA_TEMPR40[32] , 
        \R_DATA_TEMPR40[31] , \R_DATA_TEMPR40[30] , 
        \R_DATA_TEMPR40[29] , \R_DATA_TEMPR40[28] , 
        \R_DATA_TEMPR40[27] , \R_DATA_TEMPR40[26] , 
        \R_DATA_TEMPR40[25] , \R_DATA_TEMPR40[24] , 
        \R_DATA_TEMPR40[23] , \R_DATA_TEMPR40[22] , 
        \R_DATA_TEMPR40[21] , \R_DATA_TEMPR40[20] }), .B_DOUT({
        \R_DATA_TEMPR40[19] , \R_DATA_TEMPR40[18] , 
        \R_DATA_TEMPR40[17] , \R_DATA_TEMPR40[16] , 
        \R_DATA_TEMPR40[15] , \R_DATA_TEMPR40[14] , 
        \R_DATA_TEMPR40[13] , \R_DATA_TEMPR40[12] , 
        \R_DATA_TEMPR40[11] , \R_DATA_TEMPR40[10] , 
        \R_DATA_TEMPR40[9] , \R_DATA_TEMPR40[8] , \R_DATA_TEMPR40[7] , 
        \R_DATA_TEMPR40[6] , \R_DATA_TEMPR40[5] , \R_DATA_TEMPR40[4] , 
        \R_DATA_TEMPR40[3] , \R_DATA_TEMPR40[2] , \R_DATA_TEMPR40[1] , 
        \R_DATA_TEMPR40[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[40][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[10] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[10] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1422 (.A(\R_DATA_TEMPR80[3] ), .B(\R_DATA_TEMPR81[3] ), .C(
        \R_DATA_TEMPR82[3] ), .D(\R_DATA_TEMPR83[3] ), .Y(OR4_1422_Y));
    OR4 OR4_78 (.A(\R_DATA_TEMPR96[0] ), .B(\R_DATA_TEMPR97[0] ), .C(
        \R_DATA_TEMPR98[0] ), .D(\R_DATA_TEMPR99[0] ), .Y(OR4_78_Y));
    OR4 OR4_1038 (.A(OR4_1347_Y), .B(OR4_670_Y), .C(OR4_1005_Y), .D(
        OR4_196_Y), .Y(OR4_1038_Y));
    OR4 OR4_1219 (.A(OR4_948_Y), .B(OR4_1206_Y), .C(OR4_1410_Y), .D(
        OR4_1035_Y), .Y(OR4_1219_Y));
    OR4 \OR4_R_DATA[8]  (.A(OR4_818_Y), .B(OR4_1002_Y), .C(OR4_608_Y), 
        .D(OR4_1219_Y), .Y(R_DATA[8]));
    OR4 OR4_1547 (.A(\R_DATA_TEMPR112[35] ), .B(\R_DATA_TEMPR113[35] ), 
        .C(\R_DATA_TEMPR114[35] ), .D(\R_DATA_TEMPR115[35] ), .Y(
        OR4_1547_Y));
    OR4 OR4_808 (.A(\R_DATA_TEMPR116[32] ), .B(\R_DATA_TEMPR117[32] ), 
        .C(\R_DATA_TEMPR118[32] ), .D(\R_DATA_TEMPR119[32] ), .Y(
        OR4_808_Y));
    OR4 OR4_1162 (.A(\R_DATA_TEMPR96[8] ), .B(\R_DATA_TEMPR97[8] ), .C(
        \R_DATA_TEMPR98[8] ), .D(\R_DATA_TEMPR99[8] ), .Y(OR4_1162_Y));
    OR4 OR4_564 (.A(\R_DATA_TEMPR124[9] ), .B(\R_DATA_TEMPR125[9] ), 
        .C(\R_DATA_TEMPR126[9] ), .D(\R_DATA_TEMPR127[9] ), .Y(
        OR4_564_Y));
    OR4 OR4_1342 (.A(OR4_1205_Y), .B(OR4_864_Y), .C(OR4_1221_Y), .D(
        OR4_348_Y), .Y(OR4_1342_Y));
    OR4 OR4_1450 (.A(OR4_1436_Y), .B(OR4_754_Y), .C(OR4_1293_Y), .D(
        OR4_108_Y), .Y(OR4_1450_Y));
    OR4 OR4_154 (.A(\R_DATA_TEMPR4[38] ), .B(\R_DATA_TEMPR5[38] ), .C(
        \R_DATA_TEMPR6[38] ), .D(\R_DATA_TEMPR7[38] ), .Y(OR4_154_Y));
    OR2 OR2_21 (.A(\R_DATA_TEMPR84[5] ), .B(\R_DATA_TEMPR85[5] ), .Y(
        OR2_21_Y));
    OR4 OR4_727 (.A(OR4_1101_Y), .B(OR4_1364_Y), .C(OR4_870_Y), .D(
        OR4_606_Y), .Y(OR4_727_Y));
    OR4 OR4_684 (.A(\R_DATA_TEMPR40[37] ), .B(\R_DATA_TEMPR41[37] ), 
        .C(\R_DATA_TEMPR42[37] ), .D(\R_DATA_TEMPR43[37] ), .Y(
        OR4_684_Y));
    OR4 OR4_1242 (.A(OR4_1015_Y), .B(OR4_1284_Y), .C(OR4_1487_Y), .D(
        OR4_854_Y), .Y(OR4_1242_Y));
    OR4 OR4_1100 (.A(\R_DATA_TEMPR104[33] ), .B(\R_DATA_TEMPR105[33] ), 
        .C(\R_DATA_TEMPR106[33] ), .D(\R_DATA_TEMPR107[33] ), .Y(
        OR4_1100_Y));
    OR4 OR4_949 (.A(\R_DATA_TEMPR16[21] ), .B(\R_DATA_TEMPR17[21] ), 
        .C(\R_DATA_TEMPR18[21] ), .D(\R_DATA_TEMPR19[21] ), .Y(
        OR4_949_Y));
    OR4 OR4_940 (.A(OR4_324_Y), .B(OR4_589_Y), .C(OR4_571_Y), .D(
        OR4_246_Y), .Y(OR4_940_Y));
    OR4 OR4_962 (.A(OR4_799_Y), .B(OR4_626_Y), .C(OR4_19_Y), .D(
        OR4_554_Y), .Y(OR4_962_Y));
    OR4 OR4_724 (.A(OR4_860_Y), .B(OR4_117_Y), .C(OR4_758_Y), .D(
        OR4_1532_Y), .Y(OR4_724_Y));
    OR4 OR4_638 (.A(\R_DATA_TEMPR20[36] ), .B(\R_DATA_TEMPR21[36] ), 
        .C(\R_DATA_TEMPR22[36] ), .D(\R_DATA_TEMPR23[36] ), .Y(
        OR4_638_Y));
    OR4 OR4_997 (.A(\R_DATA_TEMPR100[19] ), .B(\R_DATA_TEMPR101[19] ), 
        .C(\R_DATA_TEMPR102[19] ), .D(\R_DATA_TEMPR103[19] ), .Y(
        OR4_997_Y));
    OR4 OR4_878 (.A(\R_DATA_TEMPR116[27] ), .B(\R_DATA_TEMPR117[27] ), 
        .C(\R_DATA_TEMPR118[27] ), .D(\R_DATA_TEMPR119[27] ), .Y(
        OR4_878_Y));
    OR4 OR4_1532 (.A(OR4_790_Y), .B(OR4_620_Y), .C(OR4_13_Y), .D(
        OR4_545_Y), .Y(OR4_1532_Y));
    OR4 OR4_22 (.A(\R_DATA_TEMPR16[31] ), .B(\R_DATA_TEMPR17[31] ), .C(
        \R_DATA_TEMPR18[31] ), .D(\R_DATA_TEMPR19[31] ), .Y(OR4_22_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%127%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R127C0 (.A_DOUT({
        \R_DATA_TEMPR127[39] , \R_DATA_TEMPR127[38] , 
        \R_DATA_TEMPR127[37] , \R_DATA_TEMPR127[36] , 
        \R_DATA_TEMPR127[35] , \R_DATA_TEMPR127[34] , 
        \R_DATA_TEMPR127[33] , \R_DATA_TEMPR127[32] , 
        \R_DATA_TEMPR127[31] , \R_DATA_TEMPR127[30] , 
        \R_DATA_TEMPR127[29] , \R_DATA_TEMPR127[28] , 
        \R_DATA_TEMPR127[27] , \R_DATA_TEMPR127[26] , 
        \R_DATA_TEMPR127[25] , \R_DATA_TEMPR127[24] , 
        \R_DATA_TEMPR127[23] , \R_DATA_TEMPR127[22] , 
        \R_DATA_TEMPR127[21] , \R_DATA_TEMPR127[20] }), .B_DOUT({
        \R_DATA_TEMPR127[19] , \R_DATA_TEMPR127[18] , 
        \R_DATA_TEMPR127[17] , \R_DATA_TEMPR127[16] , 
        \R_DATA_TEMPR127[15] , \R_DATA_TEMPR127[14] , 
        \R_DATA_TEMPR127[13] , \R_DATA_TEMPR127[12] , 
        \R_DATA_TEMPR127[11] , \R_DATA_TEMPR127[10] , 
        \R_DATA_TEMPR127[9] , \R_DATA_TEMPR127[8] , 
        \R_DATA_TEMPR127[7] , \R_DATA_TEMPR127[6] , 
        \R_DATA_TEMPR127[5] , \R_DATA_TEMPR127[4] , 
        \R_DATA_TEMPR127[3] , \R_DATA_TEMPR127[2] , 
        \R_DATA_TEMPR127[1] , \R_DATA_TEMPR127[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[127][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[31] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[31] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[15]  (.A(CFG3_21_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[15] ));
    OR4 OR4_1151 (.A(\R_DATA_TEMPR64[0] ), .B(\R_DATA_TEMPR65[0] ), .C(
        \R_DATA_TEMPR66[0] ), .D(\R_DATA_TEMPR67[0] ), .Y(OR4_1151_Y));
    OR4 OR4_143 (.A(OR4_478_Y), .B(OR4_1110_Y), .C(OR4_11_Y), .D(
        OR4_473_Y), .Y(OR4_143_Y));
    OR4 OR4_1444 (.A(OR4_488_Y), .B(OR4_154_Y), .C(OR4_594_Y), .D(
        OR4_417_Y), .Y(OR4_1444_Y));
    OR4 OR4_953 (.A(OR4_1569_Y), .B(OR4_242_Y), .C(OR4_1193_Y), .D(
        OR4_1004_Y), .Y(OR4_953_Y));
    OR4 OR4_632 (.A(\R_DATA_TEMPR20[24] ), .B(\R_DATA_TEMPR21[24] ), 
        .C(\R_DATA_TEMPR22[24] ), .D(\R_DATA_TEMPR23[24] ), .Y(
        OR4_632_Y));
    OR4 OR4_213 (.A(\R_DATA_TEMPR12[32] ), .B(\R_DATA_TEMPR13[32] ), 
        .C(\R_DATA_TEMPR14[32] ), .D(\R_DATA_TEMPR15[32] ), .Y(
        OR4_213_Y));
    OR4 OR4_1074 (.A(\R_DATA_TEMPR64[9] ), .B(\R_DATA_TEMPR65[9] ), .C(
        \R_DATA_TEMPR66[9] ), .D(\R_DATA_TEMPR67[9] ), .Y(OR4_1074_Y));
    OR4 OR4_821 (.A(OR4_1010_Y), .B(OR4_1400_Y), .C(OR4_1374_Y), .D(
        OR4_1037_Y), .Y(OR4_821_Y));
    OR4 OR4_201 (.A(\R_DATA_TEMPR72[21] ), .B(\R_DATA_TEMPR73[21] ), 
        .C(\R_DATA_TEMPR74[21] ), .D(\R_DATA_TEMPR75[21] ), .Y(
        OR4_201_Y));
    OR4 OR4_361 (.A(\R_DATA_TEMPR20[8] ), .B(\R_DATA_TEMPR21[8] ), .C(
        \R_DATA_TEMPR22[8] ), .D(\R_DATA_TEMPR23[8] ), .Y(OR4_361_Y));
    OR4 OR4_1244 (.A(\R_DATA_TEMPR56[2] ), .B(\R_DATA_TEMPR57[2] ), .C(
        \R_DATA_TEMPR58[2] ), .D(\R_DATA_TEMPR59[2] ), .Y(OR4_1244_Y));
    OR4 OR4_1556 (.A(\R_DATA_TEMPR28[6] ), .B(\R_DATA_TEMPR29[6] ), .C(
        \R_DATA_TEMPR30[6] ), .D(\R_DATA_TEMPR31[6] ), .Y(OR4_1556_Y));
    OR4 OR4_1373 (.A(\R_DATA_TEMPR72[39] ), .B(\R_DATA_TEMPR73[39] ), 
        .C(\R_DATA_TEMPR74[39] ), .D(\R_DATA_TEMPR75[39] ), .Y(
        OR4_1373_Y));
    OR4 OR4_856 (.A(\R_DATA_TEMPR64[3] ), .B(\R_DATA_TEMPR65[3] ), .C(
        \R_DATA_TEMPR66[3] ), .D(\R_DATA_TEMPR67[3] ), .Y(OR4_856_Y));
    OR4 OR4_751 (.A(\R_DATA_TEMPR124[19] ), .B(\R_DATA_TEMPR125[19] ), 
        .C(\R_DATA_TEMPR126[19] ), .D(\R_DATA_TEMPR127[19] ), .Y(
        OR4_751_Y));
    OR2 OR2_13 (.A(\R_DATA_TEMPR84[18] ), .B(\R_DATA_TEMPR85[18] ), .Y(
        OR2_13_Y));
    OR4 OR4_6 (.A(\R_DATA_TEMPR116[11] ), .B(\R_DATA_TEMPR117[11] ), 
        .C(\R_DATA_TEMPR118[11] ), .D(\R_DATA_TEMPR119[11] ), .Y(
        OR4_6_Y));
    OR4 OR4_918 (.A(\R_DATA_TEMPR16[2] ), .B(\R_DATA_TEMPR17[2] ), .C(
        \R_DATA_TEMPR18[2] ), .D(\R_DATA_TEMPR19[2] ), .Y(OR4_918_Y));
    OR4 OR4_1347 (.A(OR4_1147_Y), .B(OR4_560_Y), .C(OR4_793_Y), .D(
        OR4_1386_Y), .Y(OR4_1347_Y));
    OR4 OR4_271 (.A(\R_DATA_TEMPR8[0] ), .B(\R_DATA_TEMPR9[0] ), .C(
        \R_DATA_TEMPR10[0] ), .D(\R_DATA_TEMPR11[0] ), .Y(OR4_271_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%14%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C0 (.A_DOUT({
        \R_DATA_TEMPR14[39] , \R_DATA_TEMPR14[38] , 
        \R_DATA_TEMPR14[37] , \R_DATA_TEMPR14[36] , 
        \R_DATA_TEMPR14[35] , \R_DATA_TEMPR14[34] , 
        \R_DATA_TEMPR14[33] , \R_DATA_TEMPR14[32] , 
        \R_DATA_TEMPR14[31] , \R_DATA_TEMPR14[30] , 
        \R_DATA_TEMPR14[29] , \R_DATA_TEMPR14[28] , 
        \R_DATA_TEMPR14[27] , \R_DATA_TEMPR14[26] , 
        \R_DATA_TEMPR14[25] , \R_DATA_TEMPR14[24] , 
        \R_DATA_TEMPR14[23] , \R_DATA_TEMPR14[22] , 
        \R_DATA_TEMPR14[21] , \R_DATA_TEMPR14[20] }), .B_DOUT({
        \R_DATA_TEMPR14[19] , \R_DATA_TEMPR14[18] , 
        \R_DATA_TEMPR14[17] , \R_DATA_TEMPR14[16] , 
        \R_DATA_TEMPR14[15] , \R_DATA_TEMPR14[14] , 
        \R_DATA_TEMPR14[13] , \R_DATA_TEMPR14[12] , 
        \R_DATA_TEMPR14[11] , \R_DATA_TEMPR14[10] , 
        \R_DATA_TEMPR14[9] , \R_DATA_TEMPR14[8] , \R_DATA_TEMPR14[7] , 
        \R_DATA_TEMPR14[6] , \R_DATA_TEMPR14[5] , \R_DATA_TEMPR14[4] , 
        \R_DATA_TEMPR14[3] , \R_DATA_TEMPR14[2] , \R_DATA_TEMPR14[1] , 
        \R_DATA_TEMPR14[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1180 (.A(OR4_698_Y), .B(OR4_1099_Y), .C(OR4_1062_Y), .D(
        OR4_221_Y), .Y(OR4_1180_Y));
    OR4 OR4_460 (.A(\R_DATA_TEMPR116[28] ), .B(\R_DATA_TEMPR117[28] ), 
        .C(\R_DATA_TEMPR118[28] ), .D(\R_DATA_TEMPR119[28] ), .Y(
        OR4_460_Y));
    OR4 OR4_1300 (.A(\R_DATA_TEMPR44[11] ), .B(\R_DATA_TEMPR45[11] ), 
        .C(\R_DATA_TEMPR46[11] ), .D(\R_DATA_TEMPR47[11] ), .Y(
        OR4_1300_Y));
    OR4 OR4_1028 (.A(\R_DATA_TEMPR124[21] ), .B(\R_DATA_TEMPR125[21] ), 
        .C(\R_DATA_TEMPR126[21] ), .D(\R_DATA_TEMPR127[21] ), .Y(
        OR4_1028_Y));
    OR4 OR4_502 (.A(\R_DATA_TEMPR104[6] ), .B(\R_DATA_TEMPR105[6] ), 
        .C(\R_DATA_TEMPR106[6] ), .D(\R_DATA_TEMPR107[6] ), .Y(
        OR4_502_Y));
    OR4 OR4_556 (.A(OR4_1320_Y), .B(OR4_808_Y), .C(OR4_867_Y), .D(
        OR4_315_Y), .Y(OR4_556_Y));
    OR4 OR4_495 (.A(\R_DATA_TEMPR32[0] ), .B(\R_DATA_TEMPR33[0] ), .C(
        \R_DATA_TEMPR34[0] ), .D(\R_DATA_TEMPR35[0] ), .Y(OR4_495_Y));
    OR4 OR4_1192 (.A(\R_DATA_TEMPR60[27] ), .B(\R_DATA_TEMPR61[27] ), 
        .C(\R_DATA_TEMPR62[27] ), .D(\R_DATA_TEMPR63[27] ), .Y(
        OR4_1192_Y));
    OR4 OR4_1457 (.A(\R_DATA_TEMPR104[30] ), .B(\R_DATA_TEMPR105[30] ), 
        .C(\R_DATA_TEMPR106[30] ), .D(\R_DATA_TEMPR107[30] ), .Y(
        OR4_1457_Y));
    OR4 OR4_835 (.A(OR4_652_Y), .B(OR4_466_Y), .C(OR4_99_Y), .D(
        OR4_1565_Y), .Y(OR4_835_Y));
    OR4 OR4_572 (.A(OR4_1478_Y), .B(OR4_964_Y), .C(OR4_1008_Y), .D(
        OR4_874_Y), .Y(OR4_572_Y));
    OR4 OR4_618 (.A(\R_DATA_TEMPR4[39] ), .B(\R_DATA_TEMPR5[39] ), .C(
        \R_DATA_TEMPR6[39] ), .D(\R_DATA_TEMPR7[39] ), .Y(OR4_618_Y));
    OR4 OR4_1522 (.A(\R_DATA_TEMPR72[9] ), .B(\R_DATA_TEMPR73[9] ), .C(
        \R_DATA_TEMPR74[9] ), .D(\R_DATA_TEMPR75[9] ), .Y(OR4_1522_Y));
    OR4 OR4_1055 (.A(\R_DATA_TEMPR72[20] ), .B(\R_DATA_TEMPR73[20] ), 
        .C(\R_DATA_TEMPR74[20] ), .D(\R_DATA_TEMPR75[20] ), .Y(
        OR4_1055_Y));
    OR4 OR4_1037 (.A(\R_DATA_TEMPR44[38] ), .B(\R_DATA_TEMPR45[38] ), 
        .C(\R_DATA_TEMPR46[38] ), .D(\R_DATA_TEMPR47[38] ), .Y(
        OR4_1037_Y));
    CFG3 #( .INIT(8'h10) )  CFG3_8 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_8_Y));
    OR4 OR4_840 (.A(\R_DATA_TEMPR80[28] ), .B(\R_DATA_TEMPR81[28] ), 
        .C(\R_DATA_TEMPR82[28] ), .D(\R_DATA_TEMPR83[28] ), .Y(
        OR4_840_Y));
    OR4 OR4_927 (.A(\R_DATA_TEMPR4[0] ), .B(\R_DATA_TEMPR5[0] ), .C(
        \R_DATA_TEMPR6[0] ), .D(\R_DATA_TEMPR7[0] ), .Y(OR4_927_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[0]  (.A(CFG3_16_Y), .B(CFG3_2_Y)
        , .Y(\BLKY2[0] ));
    OR4 \OR4_R_DATA[17]  (.A(OR4_360_Y), .B(OR4_1124_Y), .C(OR4_1544_Y)
        , .D(OR4_66_Y), .Y(R_DATA[17]));
    OR4 OR4_142 (.A(\R_DATA_TEMPR52[27] ), .B(\R_DATA_TEMPR53[27] ), 
        .C(\R_DATA_TEMPR54[27] ), .D(\R_DATA_TEMPR55[27] ), .Y(
        OR4_142_Y));
    OR4 OR4_612 (.A(\R_DATA_TEMPR28[34] ), .B(\R_DATA_TEMPR29[34] ), 
        .C(\R_DATA_TEMPR30[34] ), .D(\R_DATA_TEMPR31[34] ), .Y(
        OR4_612_Y));
    OR4 OR4_504 (.A(\R_DATA_TEMPR72[30] ), .B(\R_DATA_TEMPR73[30] ), 
        .C(\R_DATA_TEMPR74[30] ), .D(\R_DATA_TEMPR75[30] ), .Y(
        OR4_504_Y));
    OR4 OR4_1380 (.A(\R_DATA_TEMPR12[27] ), .B(\R_DATA_TEMPR13[27] ), 
        .C(\R_DATA_TEMPR14[27] ), .D(\R_DATA_TEMPR15[27] ), .Y(
        OR4_1380_Y));
    OR4 OR4_1445 (.A(\R_DATA_TEMPR80[1] ), .B(\R_DATA_TEMPR81[1] ), .C(
        \R_DATA_TEMPR82[1] ), .D(\R_DATA_TEMPR83[1] ), .Y(OR4_1445_Y));
    OR4 OR4_945 (.A(\R_DATA_TEMPR104[24] ), .B(\R_DATA_TEMPR105[24] ), 
        .C(\R_DATA_TEMPR106[24] ), .D(\R_DATA_TEMPR107[24] ), .Y(
        OR4_945_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%71%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R71C0 (.A_DOUT({
        \R_DATA_TEMPR71[39] , \R_DATA_TEMPR71[38] , 
        \R_DATA_TEMPR71[37] , \R_DATA_TEMPR71[36] , 
        \R_DATA_TEMPR71[35] , \R_DATA_TEMPR71[34] , 
        \R_DATA_TEMPR71[33] , \R_DATA_TEMPR71[32] , 
        \R_DATA_TEMPR71[31] , \R_DATA_TEMPR71[30] , 
        \R_DATA_TEMPR71[29] , \R_DATA_TEMPR71[28] , 
        \R_DATA_TEMPR71[27] , \R_DATA_TEMPR71[26] , 
        \R_DATA_TEMPR71[25] , \R_DATA_TEMPR71[24] , 
        \R_DATA_TEMPR71[23] , \R_DATA_TEMPR71[22] , 
        \R_DATA_TEMPR71[21] , \R_DATA_TEMPR71[20] }), .B_DOUT({
        \R_DATA_TEMPR71[19] , \R_DATA_TEMPR71[18] , 
        \R_DATA_TEMPR71[17] , \R_DATA_TEMPR71[16] , 
        \R_DATA_TEMPR71[15] , \R_DATA_TEMPR71[14] , 
        \R_DATA_TEMPR71[13] , \R_DATA_TEMPR71[12] , 
        \R_DATA_TEMPR71[11] , \R_DATA_TEMPR71[10] , 
        \R_DATA_TEMPR71[9] , \R_DATA_TEMPR71[8] , \R_DATA_TEMPR71[7] , 
        \R_DATA_TEMPR71[6] , \R_DATA_TEMPR71[5] , \R_DATA_TEMPR71[4] , 
        \R_DATA_TEMPR71[3] , \R_DATA_TEMPR71[2] , \R_DATA_TEMPR71[1] , 
        \R_DATA_TEMPR71[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[71][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[17] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[17] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_902 (.A(\R_DATA_TEMPR8[36] ), .B(\R_DATA_TEMPR9[36] ), .C(
        \R_DATA_TEMPR10[36] ), .D(\R_DATA_TEMPR11[36] ), .Y(OR4_902_Y));
    OR4 OR4_1076 (.A(\R_DATA_TEMPR36[5] ), .B(\R_DATA_TEMPR37[5] ), .C(
        \R_DATA_TEMPR38[5] ), .D(\R_DATA_TEMPR39[5] ), .Y(OR4_1076_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[17]  (.A(CFG3_8_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[17] ));
    OR4 OR4_574 (.A(\R_DATA_TEMPR48[22] ), .B(\R_DATA_TEMPR49[22] ), 
        .C(\R_DATA_TEMPR50[22] ), .D(\R_DATA_TEMPR51[22] ), .Y(
        OR4_574_Y));
    OR2 OR2_11 (.A(\R_DATA_TEMPR84[21] ), .B(\R_DATA_TEMPR85[21] ), .Y(
        OR2_11_Y));
    OR4 OR4_1205 (.A(OR4_634_Y), .B(OR4_1427_Y), .C(OR4_250_Y), .D(
        OR4_566_Y), .Y(OR4_1205_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%58%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R58C0 (.A_DOUT({
        \R_DATA_TEMPR58[39] , \R_DATA_TEMPR58[38] , 
        \R_DATA_TEMPR58[37] , \R_DATA_TEMPR58[36] , 
        \R_DATA_TEMPR58[35] , \R_DATA_TEMPR58[34] , 
        \R_DATA_TEMPR58[33] , \R_DATA_TEMPR58[32] , 
        \R_DATA_TEMPR58[31] , \R_DATA_TEMPR58[30] , 
        \R_DATA_TEMPR58[29] , \R_DATA_TEMPR58[28] , 
        \R_DATA_TEMPR58[27] , \R_DATA_TEMPR58[26] , 
        \R_DATA_TEMPR58[25] , \R_DATA_TEMPR58[24] , 
        \R_DATA_TEMPR58[23] , \R_DATA_TEMPR58[22] , 
        \R_DATA_TEMPR58[21] , \R_DATA_TEMPR58[20] }), .B_DOUT({
        \R_DATA_TEMPR58[19] , \R_DATA_TEMPR58[18] , 
        \R_DATA_TEMPR58[17] , \R_DATA_TEMPR58[16] , 
        \R_DATA_TEMPR58[15] , \R_DATA_TEMPR58[14] , 
        \R_DATA_TEMPR58[13] , \R_DATA_TEMPR58[12] , 
        \R_DATA_TEMPR58[11] , \R_DATA_TEMPR58[10] , 
        \R_DATA_TEMPR58[9] , \R_DATA_TEMPR58[8] , \R_DATA_TEMPR58[7] , 
        \R_DATA_TEMPR58[6] , \R_DATA_TEMPR58[5] , \R_DATA_TEMPR58[4] , 
        \R_DATA_TEMPR58[3] , \R_DATA_TEMPR58[2] , \R_DATA_TEMPR58[1] , 
        \R_DATA_TEMPR58[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[58][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[14] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[14] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_494 (.A(\R_DATA_TEMPR0[11] ), .B(\R_DATA_TEMPR1[11] ), .C(
        \R_DATA_TEMPR2[11] ), .D(\R_DATA_TEMPR3[11] ), .Y(OR4_494_Y));
    OR4 OR4_1213 (.A(\R_DATA_TEMPR60[38] ), .B(\R_DATA_TEMPR61[38] ), 
        .C(\R_DATA_TEMPR62[38] ), .D(\R_DATA_TEMPR63[38] ), .Y(
        OR4_1213_Y));
    OR4 OR4_972 (.A(\R_DATA_TEMPR92[39] ), .B(\R_DATA_TEMPR93[39] ), 
        .C(\R_DATA_TEMPR94[39] ), .D(\R_DATA_TEMPR95[39] ), .Y(
        OR4_972_Y));
    OR4 OR4_1501 (.A(\R_DATA_TEMPR36[12] ), .B(\R_DATA_TEMPR37[12] ), 
        .C(\R_DATA_TEMPR38[12] ), .D(\R_DATA_TEMPR39[12] ), .Y(
        OR4_1501_Y));
    OR4 OR4_558 (.A(\R_DATA_TEMPR4[27] ), .B(\R_DATA_TEMPR5[27] ), .C(
        \R_DATA_TEMPR6[27] ), .D(\R_DATA_TEMPR7[27] ), .Y(OR4_558_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%81%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R81C0 (.A_DOUT({
        \R_DATA_TEMPR81[39] , \R_DATA_TEMPR81[38] , 
        \R_DATA_TEMPR81[37] , \R_DATA_TEMPR81[36] , 
        \R_DATA_TEMPR81[35] , \R_DATA_TEMPR81[34] , 
        \R_DATA_TEMPR81[33] , \R_DATA_TEMPR81[32] , 
        \R_DATA_TEMPR81[31] , \R_DATA_TEMPR81[30] , 
        \R_DATA_TEMPR81[29] , \R_DATA_TEMPR81[28] , 
        \R_DATA_TEMPR81[27] , \R_DATA_TEMPR81[26] , 
        \R_DATA_TEMPR81[25] , \R_DATA_TEMPR81[24] , 
        \R_DATA_TEMPR81[23] , \R_DATA_TEMPR81[22] , 
        \R_DATA_TEMPR81[21] , \R_DATA_TEMPR81[20] }), .B_DOUT({
        \R_DATA_TEMPR81[19] , \R_DATA_TEMPR81[18] , 
        \R_DATA_TEMPR81[17] , \R_DATA_TEMPR81[16] , 
        \R_DATA_TEMPR81[15] , \R_DATA_TEMPR81[14] , 
        \R_DATA_TEMPR81[13] , \R_DATA_TEMPR81[12] , 
        \R_DATA_TEMPR81[11] , \R_DATA_TEMPR81[10] , 
        \R_DATA_TEMPR81[9] , \R_DATA_TEMPR81[8] , \R_DATA_TEMPR81[7] , 
        \R_DATA_TEMPR81[6] , \R_DATA_TEMPR81[5] , \R_DATA_TEMPR81[4] , 
        \R_DATA_TEMPR81[3] , \R_DATA_TEMPR81[2] , \R_DATA_TEMPR81[1] , 
        \R_DATA_TEMPR81[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[81][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[20] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[20] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_55 (.A(OR4_503_Y), .B(OR4_237_Y), .C(OR4_1586_Y), .D(
        OR4_1184_Y), .Y(OR4_55_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%1%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C0 (.A_DOUT({
        \R_DATA_TEMPR1[39] , \R_DATA_TEMPR1[38] , \R_DATA_TEMPR1[37] , 
        \R_DATA_TEMPR1[36] , \R_DATA_TEMPR1[35] , \R_DATA_TEMPR1[34] , 
        \R_DATA_TEMPR1[33] , \R_DATA_TEMPR1[32] , \R_DATA_TEMPR1[31] , 
        \R_DATA_TEMPR1[30] , \R_DATA_TEMPR1[29] , \R_DATA_TEMPR1[28] , 
        \R_DATA_TEMPR1[27] , \R_DATA_TEMPR1[26] , \R_DATA_TEMPR1[25] , 
        \R_DATA_TEMPR1[24] , \R_DATA_TEMPR1[23] , \R_DATA_TEMPR1[22] , 
        \R_DATA_TEMPR1[21] , \R_DATA_TEMPR1[20] }), .B_DOUT({
        \R_DATA_TEMPR1[19] , \R_DATA_TEMPR1[18] , \R_DATA_TEMPR1[17] , 
        \R_DATA_TEMPR1[16] , \R_DATA_TEMPR1[15] , \R_DATA_TEMPR1[14] , 
        \R_DATA_TEMPR1[13] , \R_DATA_TEMPR1[12] , \R_DATA_TEMPR1[11] , 
        \R_DATA_TEMPR1[10] , \R_DATA_TEMPR1[9] , \R_DATA_TEMPR1[8] , 
        \R_DATA_TEMPR1[7] , \R_DATA_TEMPR1[6] , \R_DATA_TEMPR1[5] , 
        \R_DATA_TEMPR1[4] , \R_DATA_TEMPR1[3] , \R_DATA_TEMPR1[2] , 
        \R_DATA_TEMPR1[1] , \R_DATA_TEMPR1[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[1][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%48%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R48C0 (.A_DOUT({
        \R_DATA_TEMPR48[39] , \R_DATA_TEMPR48[38] , 
        \R_DATA_TEMPR48[37] , \R_DATA_TEMPR48[36] , 
        \R_DATA_TEMPR48[35] , \R_DATA_TEMPR48[34] , 
        \R_DATA_TEMPR48[33] , \R_DATA_TEMPR48[32] , 
        \R_DATA_TEMPR48[31] , \R_DATA_TEMPR48[30] , 
        \R_DATA_TEMPR48[29] , \R_DATA_TEMPR48[28] , 
        \R_DATA_TEMPR48[27] , \R_DATA_TEMPR48[26] , 
        \R_DATA_TEMPR48[25] , \R_DATA_TEMPR48[24] , 
        \R_DATA_TEMPR48[23] , \R_DATA_TEMPR48[22] , 
        \R_DATA_TEMPR48[21] , \R_DATA_TEMPR48[20] }), .B_DOUT({
        \R_DATA_TEMPR48[19] , \R_DATA_TEMPR48[18] , 
        \R_DATA_TEMPR48[17] , \R_DATA_TEMPR48[16] , 
        \R_DATA_TEMPR48[15] , \R_DATA_TEMPR48[14] , 
        \R_DATA_TEMPR48[13] , \R_DATA_TEMPR48[12] , 
        \R_DATA_TEMPR48[11] , \R_DATA_TEMPR48[10] , 
        \R_DATA_TEMPR48[9] , \R_DATA_TEMPR48[8] , \R_DATA_TEMPR48[7] , 
        \R_DATA_TEMPR48[6] , \R_DATA_TEMPR48[5] , \R_DATA_TEMPR48[4] , 
        \R_DATA_TEMPR48[3] , \R_DATA_TEMPR48[2] , \R_DATA_TEMPR48[1] , 
        \R_DATA_TEMPR48[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[48][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[12] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[12] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_369 (.A(\R_DATA_TEMPR76[19] ), .B(\R_DATA_TEMPR77[19] ), 
        .C(\R_DATA_TEMPR78[19] ), .D(\R_DATA_TEMPR79[19] ), .Y(
        OR4_369_Y));
    OR4 OR4_1371 (.A(\R_DATA_TEMPR24[23] ), .B(\R_DATA_TEMPR25[23] ), 
        .C(\R_DATA_TEMPR26[23] ), .D(\R_DATA_TEMPR27[23] ), .Y(
        OR4_1371_Y));
    OR4 OR4_301 (.A(\R_DATA_TEMPR32[19] ), .B(\R_DATA_TEMPR33[19] ), 
        .C(\R_DATA_TEMPR34[19] ), .D(\R_DATA_TEMPR35[19] ), .Y(
        OR4_301_Y));
    OR4 OR4_396 (.A(OR4_423_Y), .B(OR4_725_Y), .C(OR4_167_Y), .D(
        OR4_1017_Y), .Y(OR4_396_Y));
    OR4 OR4_1638 (.A(OR4_80_Y), .B(OR4_1517_Y), .C(OR4_1140_Y), .D(
        OR4_982_Y), .Y(OR4_1638_Y));
    OR4 OR4_249 (.A(\R_DATA_TEMPR96[33] ), .B(\R_DATA_TEMPR97[33] ), 
        .C(\R_DATA_TEMPR98[33] ), .D(\R_DATA_TEMPR99[33] ), .Y(
        OR4_249_Y));
    OR4 OR4_371 (.A(\R_DATA_TEMPR60[0] ), .B(\R_DATA_TEMPR61[0] ), .C(
        \R_DATA_TEMPR62[0] ), .D(\R_DATA_TEMPR63[0] ), .Y(OR4_371_Y));
    OR4 OR4_425 (.A(\R_DATA_TEMPR44[0] ), .B(\R_DATA_TEMPR45[0] ), .C(
        \R_DATA_TEMPR46[0] ), .D(\R_DATA_TEMPR47[0] ), .Y(OR4_425_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%10%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C0 (.A_DOUT({
        \R_DATA_TEMPR10[39] , \R_DATA_TEMPR10[38] , 
        \R_DATA_TEMPR10[37] , \R_DATA_TEMPR10[36] , 
        \R_DATA_TEMPR10[35] , \R_DATA_TEMPR10[34] , 
        \R_DATA_TEMPR10[33] , \R_DATA_TEMPR10[32] , 
        \R_DATA_TEMPR10[31] , \R_DATA_TEMPR10[30] , 
        \R_DATA_TEMPR10[29] , \R_DATA_TEMPR10[28] , 
        \R_DATA_TEMPR10[27] , \R_DATA_TEMPR10[26] , 
        \R_DATA_TEMPR10[25] , \R_DATA_TEMPR10[24] , 
        \R_DATA_TEMPR10[23] , \R_DATA_TEMPR10[22] , 
        \R_DATA_TEMPR10[21] , \R_DATA_TEMPR10[20] }), .B_DOUT({
        \R_DATA_TEMPR10[19] , \R_DATA_TEMPR10[18] , 
        \R_DATA_TEMPR10[17] , \R_DATA_TEMPR10[16] , 
        \R_DATA_TEMPR10[15] , \R_DATA_TEMPR10[14] , 
        \R_DATA_TEMPR10[13] , \R_DATA_TEMPR10[12] , 
        \R_DATA_TEMPR10[11] , \R_DATA_TEMPR10[10] , 
        \R_DATA_TEMPR10[9] , \R_DATA_TEMPR10[8] , \R_DATA_TEMPR10[7] , 
        \R_DATA_TEMPR10[6] , \R_DATA_TEMPR10[5] , \R_DATA_TEMPR10[4] , 
        \R_DATA_TEMPR10[3] , \R_DATA_TEMPR10[2] , \R_DATA_TEMPR10[1] , 
        \R_DATA_TEMPR10[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[2] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_815 (.A(\R_DATA_TEMPR104[25] ), .B(\R_DATA_TEMPR105[25] ), 
        .C(\R_DATA_TEMPR106[25] ), .D(\R_DATA_TEMPR107[25] ), .Y(
        OR4_815_Y));
    OR4 OR4_400 (.A(OR4_111_Y), .B(OR4_100_Y), .C(OR4_628_Y), .D(
        OR4_1082_Y), .Y(OR4_400_Y));
    OR4 OR4_1568 (.A(OR4_1379_Y), .B(OR4_1201_Y), .C(OR4_1336_Y), .D(
        OR4_1335_Y), .Y(OR4_1568_Y));
    OR4 \OR4_R_DATA[38]  (.A(OR4_314_Y), .B(OR4_85_Y), .C(OR4_962_Y), 
        .D(OR4_1187_Y), .Y(R_DATA[38]));
    OR4 OR4_636 (.A(\R_DATA_TEMPR64[33] ), .B(\R_DATA_TEMPR65[33] ), 
        .C(\R_DATA_TEMPR66[33] ), .D(\R_DATA_TEMPR67[33] ), .Y(
        OR4_636_Y));
    OR4 OR4_456 (.A(\R_DATA_TEMPR68[6] ), .B(\R_DATA_TEMPR69[6] ), .C(
        \R_DATA_TEMPR70[6] ), .D(\R_DATA_TEMPR71[6] ), .Y(OR4_456_Y));
    OR4 OR4_1027 (.A(\R_DATA_TEMPR68[23] ), .B(\R_DATA_TEMPR69[23] ), 
        .C(\R_DATA_TEMPR70[23] ), .D(\R_DATA_TEMPR71[23] ), .Y(
        OR4_1027_Y));
    OR4 OR4_1346 (.A(\R_DATA_TEMPR28[18] ), .B(\R_DATA_TEMPR29[18] ), 
        .C(\R_DATA_TEMPR30[18] ), .D(\R_DATA_TEMPR31[18] ), .Y(
        OR4_1346_Y));
    OR4 OR4_1285 (.A(\R_DATA_TEMPR104[32] ), .B(\R_DATA_TEMPR105[32] ), 
        .C(\R_DATA_TEMPR106[32] ), .D(\R_DATA_TEMPR107[32] ), .Y(
        OR4_1285_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[5]  (.A(CFG3_11_Y), .B(CFG3_2_Y)
        , .Y(\BLKY2[5] ));
    OR4 OR4_1119 (.A(OR4_1253_Y), .B(OR4_1558_Y), .C(OR4_999_Y), .D(
        OR4_232_Y), .Y(OR4_1119_Y));
    OR4 OR4_1269 (.A(\R_DATA_TEMPR116[31] ), .B(\R_DATA_TEMPR117[31] ), 
        .C(\R_DATA_TEMPR118[31] ), .D(\R_DATA_TEMPR119[31] ), .Y(
        OR4_1269_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%22%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C0 (.A_DOUT({
        \R_DATA_TEMPR22[39] , \R_DATA_TEMPR22[38] , 
        \R_DATA_TEMPR22[37] , \R_DATA_TEMPR22[36] , 
        \R_DATA_TEMPR22[35] , \R_DATA_TEMPR22[34] , 
        \R_DATA_TEMPR22[33] , \R_DATA_TEMPR22[32] , 
        \R_DATA_TEMPR22[31] , \R_DATA_TEMPR22[30] , 
        \R_DATA_TEMPR22[29] , \R_DATA_TEMPR22[28] , 
        \R_DATA_TEMPR22[27] , \R_DATA_TEMPR22[26] , 
        \R_DATA_TEMPR22[25] , \R_DATA_TEMPR22[24] , 
        \R_DATA_TEMPR22[23] , \R_DATA_TEMPR22[22] , 
        \R_DATA_TEMPR22[21] , \R_DATA_TEMPR22[20] }), .B_DOUT({
        \R_DATA_TEMPR22[19] , \R_DATA_TEMPR22[18] , 
        \R_DATA_TEMPR22[17] , \R_DATA_TEMPR22[16] , 
        \R_DATA_TEMPR22[15] , \R_DATA_TEMPR22[14] , 
        \R_DATA_TEMPR22[13] , \R_DATA_TEMPR22[12] , 
        \R_DATA_TEMPR22[11] , \R_DATA_TEMPR22[10] , 
        \R_DATA_TEMPR22[9] , \R_DATA_TEMPR22[8] , \R_DATA_TEMPR22[7] , 
        \R_DATA_TEMPR22[6] , \R_DATA_TEMPR22[5] , \R_DATA_TEMPR22[4] , 
        \R_DATA_TEMPR22[3] , \R_DATA_TEMPR22[2] , \R_DATA_TEMPR22[1] , 
        \R_DATA_TEMPR22[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%34%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R34C0 (.A_DOUT({
        \R_DATA_TEMPR34[39] , \R_DATA_TEMPR34[38] , 
        \R_DATA_TEMPR34[37] , \R_DATA_TEMPR34[36] , 
        \R_DATA_TEMPR34[35] , \R_DATA_TEMPR34[34] , 
        \R_DATA_TEMPR34[33] , \R_DATA_TEMPR34[32] , 
        \R_DATA_TEMPR34[31] , \R_DATA_TEMPR34[30] , 
        \R_DATA_TEMPR34[29] , \R_DATA_TEMPR34[28] , 
        \R_DATA_TEMPR34[27] , \R_DATA_TEMPR34[26] , 
        \R_DATA_TEMPR34[25] , \R_DATA_TEMPR34[24] , 
        \R_DATA_TEMPR34[23] , \R_DATA_TEMPR34[22] , 
        \R_DATA_TEMPR34[21] , \R_DATA_TEMPR34[20] }), .B_DOUT({
        \R_DATA_TEMPR34[19] , \R_DATA_TEMPR34[18] , 
        \R_DATA_TEMPR34[17] , \R_DATA_TEMPR34[16] , 
        \R_DATA_TEMPR34[15] , \R_DATA_TEMPR34[14] , 
        \R_DATA_TEMPR34[13] , \R_DATA_TEMPR34[12] , 
        \R_DATA_TEMPR34[11] , \R_DATA_TEMPR34[10] , 
        \R_DATA_TEMPR34[9] , \R_DATA_TEMPR34[8] , \R_DATA_TEMPR34[7] , 
        \R_DATA_TEMPR34[6] , \R_DATA_TEMPR34[5] , \R_DATA_TEMPR34[4] , 
        \R_DATA_TEMPR34[3] , \R_DATA_TEMPR34[2] , \R_DATA_TEMPR34[1] , 
        \R_DATA_TEMPR34[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[34][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[8] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[8] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_888 (.A(\R_DATA_TEMPR72[35] ), .B(\R_DATA_TEMPR73[35] ), 
        .C(\R_DATA_TEMPR74[35] ), .D(\R_DATA_TEMPR75[35] ), .Y(
        OR4_888_Y));
    OR4 OR4_470 (.A(\R_DATA_TEMPR124[24] ), .B(\R_DATA_TEMPR125[24] ), 
        .C(\R_DATA_TEMPR126[24] ), .D(\R_DATA_TEMPR127[24] ), .Y(
        OR4_470_Y));
    OR4 OR4_1581 (.A(\R_DATA_TEMPR100[20] ), .B(\R_DATA_TEMPR101[20] ), 
        .C(\R_DATA_TEMPR102[20] ), .D(\R_DATA_TEMPR103[20] ), .Y(
        OR4_1581_Y));
    OR4 OR4_849 (.A(\R_DATA_TEMPR96[22] ), .B(\R_DATA_TEMPR97[22] ), 
        .C(\R_DATA_TEMPR98[22] ), .D(\R_DATA_TEMPR99[22] ), .Y(
        OR4_849_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%115%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R115C0 (.A_DOUT({
        \R_DATA_TEMPR115[39] , \R_DATA_TEMPR115[38] , 
        \R_DATA_TEMPR115[37] , \R_DATA_TEMPR115[36] , 
        \R_DATA_TEMPR115[35] , \R_DATA_TEMPR115[34] , 
        \R_DATA_TEMPR115[33] , \R_DATA_TEMPR115[32] , 
        \R_DATA_TEMPR115[31] , \R_DATA_TEMPR115[30] , 
        \R_DATA_TEMPR115[29] , \R_DATA_TEMPR115[28] , 
        \R_DATA_TEMPR115[27] , \R_DATA_TEMPR115[26] , 
        \R_DATA_TEMPR115[25] , \R_DATA_TEMPR115[24] , 
        \R_DATA_TEMPR115[23] , \R_DATA_TEMPR115[22] , 
        \R_DATA_TEMPR115[21] , \R_DATA_TEMPR115[20] }), .B_DOUT({
        \R_DATA_TEMPR115[19] , \R_DATA_TEMPR115[18] , 
        \R_DATA_TEMPR115[17] , \R_DATA_TEMPR115[16] , 
        \R_DATA_TEMPR115[15] , \R_DATA_TEMPR115[14] , 
        \R_DATA_TEMPR115[13] , \R_DATA_TEMPR115[12] , 
        \R_DATA_TEMPR115[11] , \R_DATA_TEMPR115[10] , 
        \R_DATA_TEMPR115[9] , \R_DATA_TEMPR115[8] , 
        \R_DATA_TEMPR115[7] , \R_DATA_TEMPR115[6] , 
        \R_DATA_TEMPR115[5] , \R_DATA_TEMPR115[4] , 
        \R_DATA_TEMPR115[3] , \R_DATA_TEMPR115[2] , 
        \R_DATA_TEMPR115[1] , \R_DATA_TEMPR115[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[115][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[28] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[28] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1150 (.A(\R_DATA_TEMPR124[13] ), .B(\R_DATA_TEMPR125[13] ), 
        .C(\R_DATA_TEMPR126[13] ), .D(\R_DATA_TEMPR127[13] ), .Y(
        OR4_1150_Y));
    OR4 OR4_352 (.A(\R_DATA_TEMPR8[19] ), .B(\R_DATA_TEMPR9[19] ), .C(
        \R_DATA_TEMPR10[19] ), .D(\R_DATA_TEMPR11[19] ), .Y(OR4_352_Y));
    OR4 OR4_15 (.A(\R_DATA_TEMPR16[0] ), .B(\R_DATA_TEMPR17[0] ), .C(
        \R_DATA_TEMPR18[0] ), .D(\R_DATA_TEMPR19[0] ), .Y(OR4_15_Y));
    OR4 OR4_1606 (.A(\R_DATA_TEMPR40[0] ), .B(\R_DATA_TEMPR41[0] ), .C(
        \R_DATA_TEMPR42[0] ), .D(\R_DATA_TEMPR43[0] ), .Y(OR4_1606_Y));
    OR4 OR4_424 (.A(OR4_863_Y), .B(OR2_33_Y), .C(\R_DATA_TEMPR86[6] ), 
        .D(\R_DATA_TEMPR87[6] ), .Y(OR4_424_Y));
    OR4 OR4_281 (.A(\R_DATA_TEMPR104[12] ), .B(\R_DATA_TEMPR105[12] ), 
        .C(\R_DATA_TEMPR106[12] ), .D(\R_DATA_TEMPR107[12] ), .Y(
        OR4_281_Y));
    OR4 OR4_769 (.A(OR4_894_Y), .B(OR4_402_Y), .C(OR4_449_Y), .D(
        OR4_807_Y), .Y(OR4_769_Y));
    OR4 OR4_1635 (.A(\R_DATA_TEMPR108[27] ), .B(\R_DATA_TEMPR109[27] ), 
        .C(\R_DATA_TEMPR110[27] ), .D(\R_DATA_TEMPR111[27] ), .Y(
        OR4_1635_Y));
    OR4 OR4_1628 (.A(\R_DATA_TEMPR72[5] ), .B(\R_DATA_TEMPR73[5] ), .C(
        \R_DATA_TEMPR74[5] ), .D(\R_DATA_TEMPR75[5] ), .Y(OR4_1628_Y));
    OR4 OR4_1116 (.A(\R_DATA_TEMPR60[18] ), .B(\R_DATA_TEMPR61[18] ), 
        .C(\R_DATA_TEMPR62[18] ), .D(\R_DATA_TEMPR63[18] ), .Y(
        OR4_1116_Y));
    OR4 OR4_864 (.A(OR4_795_Y), .B(OR4_609_Y), .C(OR4_245_Y), .D(
        OR4_81_Y), .Y(OR4_864_Y));
    OR4 OR4_194 (.A(\R_DATA_TEMPR52[21] ), .B(\R_DATA_TEMPR53[21] ), 
        .C(\R_DATA_TEMPR54[21] ), .D(\R_DATA_TEMPR55[21] ), .Y(
        OR4_194_Y));
    OR4 OR4_326 (.A(OR4_1589_Y), .B(OR4_75_Y), .C(OR4_613_Y), .D(
        OR4_1_Y), .Y(OR4_326_Y));
    OR4 OR4_1411 (.A(\R_DATA_TEMPR48[5] ), .B(\R_DATA_TEMPR49[5] ), .C(
        \R_DATA_TEMPR50[5] ), .D(\R_DATA_TEMPR51[5] ), .Y(OR4_1411_Y));
    OR4 OR4_1448 (.A(OR4_633_Y), .B(OR4_1497_Y), .C(OR4_655_Y), .D(
        OR4_911_Y), .Y(OR4_1448_Y));
    OR4 OR4_1237 (.A(\R_DATA_TEMPR60[21] ), .B(\R_DATA_TEMPR61[21] ), 
        .C(\R_DATA_TEMPR62[21] ), .D(\R_DATA_TEMPR63[21] ), .Y(
        OR4_1237_Y));
    OR4 OR4_1598 (.A(\R_DATA_TEMPR112[15] ), .B(\R_DATA_TEMPR113[15] ), 
        .C(\R_DATA_TEMPR114[15] ), .D(\R_DATA_TEMPR115[15] ), .Y(
        OR4_1598_Y));
    OR4 OR4_747 (.A(\R_DATA_TEMPR36[31] ), .B(\R_DATA_TEMPR37[31] ), 
        .C(\R_DATA_TEMPR38[31] ), .D(\R_DATA_TEMPR39[31] ), .Y(
        OR4_747_Y));
    OR4 OR4_563 (.A(OR4_680_Y), .B(OR4_987_Y), .C(OR4_1233_Y), .D(
        OR4_1033_Y), .Y(OR4_563_Y));
    OR4 OR4_93 (.A(\R_DATA_TEMPR112[14] ), .B(\R_DATA_TEMPR113[14] ), 
        .C(\R_DATA_TEMPR114[14] ), .D(\R_DATA_TEMPR115[14] ), .Y(
        OR4_93_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%57%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R57C0 (.A_DOUT({
        \R_DATA_TEMPR57[39] , \R_DATA_TEMPR57[38] , 
        \R_DATA_TEMPR57[37] , \R_DATA_TEMPR57[36] , 
        \R_DATA_TEMPR57[35] , \R_DATA_TEMPR57[34] , 
        \R_DATA_TEMPR57[33] , \R_DATA_TEMPR57[32] , 
        \R_DATA_TEMPR57[31] , \R_DATA_TEMPR57[30] , 
        \R_DATA_TEMPR57[29] , \R_DATA_TEMPR57[28] , 
        \R_DATA_TEMPR57[27] , \R_DATA_TEMPR57[26] , 
        \R_DATA_TEMPR57[25] , \R_DATA_TEMPR57[24] , 
        \R_DATA_TEMPR57[23] , \R_DATA_TEMPR57[22] , 
        \R_DATA_TEMPR57[21] , \R_DATA_TEMPR57[20] }), .B_DOUT({
        \R_DATA_TEMPR57[19] , \R_DATA_TEMPR57[18] , 
        \R_DATA_TEMPR57[17] , \R_DATA_TEMPR57[16] , 
        \R_DATA_TEMPR57[15] , \R_DATA_TEMPR57[14] , 
        \R_DATA_TEMPR57[13] , \R_DATA_TEMPR57[12] , 
        \R_DATA_TEMPR57[11] , \R_DATA_TEMPR57[10] , 
        \R_DATA_TEMPR57[9] , \R_DATA_TEMPR57[8] , \R_DATA_TEMPR57[7] , 
        \R_DATA_TEMPR57[6] , \R_DATA_TEMPR57[5] , \R_DATA_TEMPR57[4] , 
        \R_DATA_TEMPR57[3] , \R_DATA_TEMPR57[2] , \R_DATA_TEMPR57[1] , 
        \R_DATA_TEMPR57[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[57][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[14] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[14] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1211 (.A(OR4_1299_Y), .B(OR4_1103_Y), .C(OR4_736_Y), .D(
        OR4_579_Y), .Y(OR4_1211_Y));
    OR4 OR4_744 (.A(\R_DATA_TEMPR8[13] ), .B(\R_DATA_TEMPR9[13] ), .C(
        \R_DATA_TEMPR10[13] ), .D(\R_DATA_TEMPR11[13] ), .Y(OR4_744_Y));
    OR4 OR4_1350 (.A(\R_DATA_TEMPR68[20] ), .B(\R_DATA_TEMPR69[20] ), 
        .C(\R_DATA_TEMPR70[20] ), .D(\R_DATA_TEMPR71[20] ), .Y(
        OR4_1350_Y));
    OR4 OR4_616 (.A(\R_DATA_TEMPR44[12] ), .B(\R_DATA_TEMPR45[12] ), 
        .C(\R_DATA_TEMPR46[12] ), .D(\R_DATA_TEMPR47[12] ), .Y(
        OR4_616_Y));
    OR4 OR4_309 (.A(\R_DATA_TEMPR120[0] ), .B(\R_DATA_TEMPR121[0] ), 
        .C(\R_DATA_TEMPR122[0] ), .D(\R_DATA_TEMPR123[0] ), .Y(
        OR4_309_Y));
    OR4 OR4_1118 (.A(\R_DATA_TEMPR112[33] ), .B(\R_DATA_TEMPR113[33] ), 
        .C(\R_DATA_TEMPR114[33] ), .D(\R_DATA_TEMPR115[33] ), .Y(
        OR4_1118_Y));
    OR4 OR4_582 (.A(\R_DATA_TEMPR60[31] ), .B(\R_DATA_TEMPR61[31] ), 
        .C(\R_DATA_TEMPR62[31] ), .D(\R_DATA_TEMPR63[31] ), .Y(
        OR4_582_Y));
    OR4 OR4_24 (.A(\R_DATA_TEMPR24[1] ), .B(\R_DATA_TEMPR25[1] ), .C(
        \R_DATA_TEMPR26[1] ), .D(\R_DATA_TEMPR27[1] ), .Y(OR4_24_Y));
    OR4 OR4_1299 (.A(\R_DATA_TEMPR16[13] ), .B(\R_DATA_TEMPR17[13] ), 
        .C(\R_DATA_TEMPR18[13] ), .D(\R_DATA_TEMPR19[13] ), .Y(
        OR4_1299_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%47%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R47C0 (.A_DOUT({
        \R_DATA_TEMPR47[39] , \R_DATA_TEMPR47[38] , 
        \R_DATA_TEMPR47[37] , \R_DATA_TEMPR47[36] , 
        \R_DATA_TEMPR47[35] , \R_DATA_TEMPR47[34] , 
        \R_DATA_TEMPR47[33] , \R_DATA_TEMPR47[32] , 
        \R_DATA_TEMPR47[31] , \R_DATA_TEMPR47[30] , 
        \R_DATA_TEMPR47[29] , \R_DATA_TEMPR47[28] , 
        \R_DATA_TEMPR47[27] , \R_DATA_TEMPR47[26] , 
        \R_DATA_TEMPR47[25] , \R_DATA_TEMPR47[24] , 
        \R_DATA_TEMPR47[23] , \R_DATA_TEMPR47[22] , 
        \R_DATA_TEMPR47[21] , \R_DATA_TEMPR47[20] }), .B_DOUT({
        \R_DATA_TEMPR47[19] , \R_DATA_TEMPR47[18] , 
        \R_DATA_TEMPR47[17] , \R_DATA_TEMPR47[16] , 
        \R_DATA_TEMPR47[15] , \R_DATA_TEMPR47[14] , 
        \R_DATA_TEMPR47[13] , \R_DATA_TEMPR47[12] , 
        \R_DATA_TEMPR47[11] , \R_DATA_TEMPR47[10] , 
        \R_DATA_TEMPR47[9] , \R_DATA_TEMPR47[8] , \R_DATA_TEMPR47[7] , 
        \R_DATA_TEMPR47[6] , \R_DATA_TEMPR47[5] , \R_DATA_TEMPR47[4] , 
        \R_DATA_TEMPR47[3] , \R_DATA_TEMPR47[2] , \R_DATA_TEMPR47[1] , 
        \R_DATA_TEMPR47[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[47][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[11] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[11] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_993 (.A(\R_DATA_TEMPR96[20] ), .B(\R_DATA_TEMPR97[20] ), 
        .C(\R_DATA_TEMPR98[20] ), .D(\R_DATA_TEMPR99[20] ), .Y(
        OR4_993_Y));
    OR4 OR4_8 (.A(OR4_1216_Y), .B(OR4_153_Y), .C(OR4_945_Y), .D(
        OR4_1202_Y), .Y(OR4_8_Y));
    OR4 OR4_1632 (.A(\R_DATA_TEMPR36[23] ), .B(\R_DATA_TEMPR37[23] ), 
        .C(\R_DATA_TEMPR38[23] ), .D(\R_DATA_TEMPR39[23] ), .Y(
        OR4_1632_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[7]  (.A(CFG3_21_Y), .B(CFG3_2_Y)
        , .Y(\BLKY2[7] ));
    OR4 OR4_379 (.A(\R_DATA_TEMPR60[5] ), .B(\R_DATA_TEMPR61[5] ), .C(
        \R_DATA_TEMPR62[5] ), .D(\R_DATA_TEMPR63[5] ), .Y(OR4_379_Y));
    OR4 OR4_1436 (.A(\R_DATA_TEMPR32[3] ), .B(\R_DATA_TEMPR33[3] ), .C(
        \R_DATA_TEMPR34[3] ), .D(\R_DATA_TEMPR35[3] ), .Y(OR4_1436_Y));
    OR4 OR4_1334 (.A(\R_DATA_TEMPR64[35] ), .B(\R_DATA_TEMPR65[35] ), 
        .C(\R_DATA_TEMPR66[35] ), .D(\R_DATA_TEMPR67[35] ), .Y(
        OR4_1334_Y));
    OR4 OR4_1004 (.A(OR4_1413_Y), .B(OR4_79_Y), .C(OR4_1146_Y), .D(
        OR4_381_Y), .Y(OR4_1004_Y));
    OR4 OR4_841 (.A(\R_DATA_TEMPR92[25] ), .B(\R_DATA_TEMPR93[25] ), 
        .C(\R_DATA_TEMPR94[25] ), .D(\R_DATA_TEMPR95[25] ), .Y(
        OR4_841_Y));
    OR4 OR4_250 (.A(\R_DATA_TEMPR8[10] ), .B(\R_DATA_TEMPR9[10] ), .C(
        \R_DATA_TEMPR10[10] ), .D(\R_DATA_TEMPR11[10] ), .Y(OR4_250_Y));
    OR4 OR4_1172 (.A(\R_DATA_TEMPR116[34] ), .B(\R_DATA_TEMPR117[34] ), 
        .C(\R_DATA_TEMPR118[34] ), .D(\R_DATA_TEMPR119[34] ), .Y(
        OR4_1172_Y));
    OR4 OR4_557 (.A(\R_DATA_TEMPR20[31] ), .B(\R_DATA_TEMPR21[31] ), 
        .C(\R_DATA_TEMPR22[31] ), .D(\R_DATA_TEMPR23[31] ), .Y(
        OR4_557_Y));
    OR4 OR4_896 (.A(\R_DATA_TEMPR120[16] ), .B(\R_DATA_TEMPR121[16] ), 
        .C(\R_DATA_TEMPR122[16] ), .D(\R_DATA_TEMPR123[16] ), .Y(
        OR4_896_Y));
    OR2 OR2_4 (.A(\R_DATA_TEMPR84[7] ), .B(\R_DATA_TEMPR85[7] ), .Y(
        OR2_4_Y));
    OR4 OR4_334 (.A(\R_DATA_TEMPR48[14] ), .B(\R_DATA_TEMPR49[14] ), 
        .C(\R_DATA_TEMPR50[14] ), .D(\R_DATA_TEMPR51[14] ), .Y(
        OR4_334_Y));
    OR4 OR4_791 (.A(\R_DATA_TEMPR8[27] ), .B(\R_DATA_TEMPR9[27] ), .C(
        \R_DATA_TEMPR10[27] ), .D(\R_DATA_TEMPR11[27] ), .Y(OR4_791_Y));
    OR4 OR4_1303 (.A(\R_DATA_TEMPR76[9] ), .B(\R_DATA_TEMPR77[9] ), .C(
        \R_DATA_TEMPR78[9] ), .D(\R_DATA_TEMPR79[9] ), .Y(OR4_1303_Y));
    OR4 OR4_1144 (.A(\R_DATA_TEMPR8[14] ), .B(\R_DATA_TEMPR9[14] ), .C(
        \R_DATA_TEMPR10[14] ), .D(\R_DATA_TEMPR11[14] ), .Y(OR4_1144_Y)
        );
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%30%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C0 (.A_DOUT({
        \R_DATA_TEMPR30[39] , \R_DATA_TEMPR30[38] , 
        \R_DATA_TEMPR30[37] , \R_DATA_TEMPR30[36] , 
        \R_DATA_TEMPR30[35] , \R_DATA_TEMPR30[34] , 
        \R_DATA_TEMPR30[33] , \R_DATA_TEMPR30[32] , 
        \R_DATA_TEMPR30[31] , \R_DATA_TEMPR30[30] , 
        \R_DATA_TEMPR30[29] , \R_DATA_TEMPR30[28] , 
        \R_DATA_TEMPR30[27] , \R_DATA_TEMPR30[26] , 
        \R_DATA_TEMPR30[25] , \R_DATA_TEMPR30[24] , 
        \R_DATA_TEMPR30[23] , \R_DATA_TEMPR30[22] , 
        \R_DATA_TEMPR30[21] , \R_DATA_TEMPR30[20] }), .B_DOUT({
        \R_DATA_TEMPR30[19] , \R_DATA_TEMPR30[18] , 
        \R_DATA_TEMPR30[17] , \R_DATA_TEMPR30[16] , 
        \R_DATA_TEMPR30[15] , \R_DATA_TEMPR30[14] , 
        \R_DATA_TEMPR30[13] , \R_DATA_TEMPR30[12] , 
        \R_DATA_TEMPR30[11] , \R_DATA_TEMPR30[10] , 
        \R_DATA_TEMPR30[9] , \R_DATA_TEMPR30[8] , \R_DATA_TEMPR30[7] , 
        \R_DATA_TEMPR30[6] , \R_DATA_TEMPR30[5] , \R_DATA_TEMPR30[4] , 
        \R_DATA_TEMPR30[3] , \R_DATA_TEMPR30[2] , \R_DATA_TEMPR30[1] , 
        \R_DATA_TEMPR30[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_131 (.A(\R_DATA_TEMPR24[36] ), .B(\R_DATA_TEMPR25[36] ), 
        .C(\R_DATA_TEMPR26[36] ), .D(\R_DATA_TEMPR27[36] ), .Y(
        OR4_131_Y));
    OR4 OR4_584 (.A(\R_DATA_TEMPR96[9] ), .B(\R_DATA_TEMPR97[9] ), .C(
        \R_DATA_TEMPR98[9] ), .D(\R_DATA_TEMPR99[9] ), .Y(OR4_584_Y));
    OR4 OR4_1637 (.A(OR4_1437_Y), .B(OR2_23_Y), .C(
        \R_DATA_TEMPR86[29] ), .D(\R_DATA_TEMPR87[29] ), .Y(OR4_1637_Y)
        );
    OR4 OR4_659 (.A(\R_DATA_TEMPR52[31] ), .B(\R_DATA_TEMPR53[31] ), 
        .C(\R_DATA_TEMPR54[31] ), .D(\R_DATA_TEMPR55[31] ), .Y(
        OR4_659_Y));
    OR4 OR4_1540 (.A(\R_DATA_TEMPR0[14] ), .B(\R_DATA_TEMPR1[14] ), .C(
        \R_DATA_TEMPR2[14] ), .D(\R_DATA_TEMPR3[14] ), .Y(OR4_1540_Y));
    OR4 OR4_982 (.A(\R_DATA_TEMPR28[14] ), .B(\R_DATA_TEMPR29[14] ), 
        .C(\R_DATA_TEMPR30[14] ), .D(\R_DATA_TEMPR31[14] ), .Y(
        OR4_982_Y));
    OR4 OR4_596 (.A(\R_DATA_TEMPR120[27] ), .B(\R_DATA_TEMPR121[27] ), 
        .C(\R_DATA_TEMPR122[27] ), .D(\R_DATA_TEMPR123[27] ), .Y(
        OR4_596_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[8]  (.A(CFG3_13_Y), .B(CFG3_4_Y)
        , .Y(\BLKX2[8] ));
    OR4 \OR4_R_DATA[39]  (.A(OR4_899_Y), .B(OR4_544_Y), .C(OR4_428_Y), 
        .D(OR4_133_Y), .Y(R_DATA[39]));
    OR4 OR4_1625 (.A(\R_DATA_TEMPR72[36] ), .B(\R_DATA_TEMPR73[36] ), 
        .C(\R_DATA_TEMPR74[36] ), .D(\R_DATA_TEMPR75[36] ), .Y(
        OR4_1625_Y));
    OR4 OR4_256 (.A(\R_DATA_TEMPR32[35] ), .B(\R_DATA_TEMPR33[35] ), 
        .C(\R_DATA_TEMPR34[35] ), .D(\R_DATA_TEMPR35[35] ), .Y(
        OR4_256_Y));
    OR2 OR2_0 (.A(\R_DATA_TEMPR84[16] ), .B(\R_DATA_TEMPR85[16] ), .Y(
        OR2_0_Y));
    OR4 OR4_1255 (.A(\R_DATA_TEMPR76[8] ), .B(\R_DATA_TEMPR77[8] ), .C(
        \R_DATA_TEMPR78[8] ), .D(\R_DATA_TEMPR79[8] ), .Y(OR4_1255_Y));
    OR4 OR4_1084 (.A(\R_DATA_TEMPR96[25] ), .B(\R_DATA_TEMPR97[25] ), 
        .C(\R_DATA_TEMPR98[25] ), .D(\R_DATA_TEMPR99[25] ), .Y(
        OR4_1084_Y));
    OR4 OR4_75 (.A(\R_DATA_TEMPR36[28] ), .B(\R_DATA_TEMPR37[28] ), .C(
        \R_DATA_TEMPR38[28] ), .D(\R_DATA_TEMPR39[28] ), .Y(OR4_75_Y));
    OR4 OR4_1248 (.A(OR4_537_Y), .B(OR4_782_Y), .C(OR4_300_Y), .D(
        OR4_25_Y), .Y(OR4_1248_Y));
    OR2 OR2_6 (.A(\R_DATA_TEMPR84[3] ), .B(\R_DATA_TEMPR85[3] ), .Y(
        OR2_6_Y));
    OR4 OR4_1339 (.A(\R_DATA_TEMPR68[9] ), .B(\R_DATA_TEMPR69[9] ), .C(
        \R_DATA_TEMPR70[9] ), .D(\R_DATA_TEMPR71[9] ), .Y(OR4_1339_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%121%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R121C0 (.A_DOUT({
        \R_DATA_TEMPR121[39] , \R_DATA_TEMPR121[38] , 
        \R_DATA_TEMPR121[37] , \R_DATA_TEMPR121[36] , 
        \R_DATA_TEMPR121[35] , \R_DATA_TEMPR121[34] , 
        \R_DATA_TEMPR121[33] , \R_DATA_TEMPR121[32] , 
        \R_DATA_TEMPR121[31] , \R_DATA_TEMPR121[30] , 
        \R_DATA_TEMPR121[29] , \R_DATA_TEMPR121[28] , 
        \R_DATA_TEMPR121[27] , \R_DATA_TEMPR121[26] , 
        \R_DATA_TEMPR121[25] , \R_DATA_TEMPR121[24] , 
        \R_DATA_TEMPR121[23] , \R_DATA_TEMPR121[22] , 
        \R_DATA_TEMPR121[21] , \R_DATA_TEMPR121[20] }), .B_DOUT({
        \R_DATA_TEMPR121[19] , \R_DATA_TEMPR121[18] , 
        \R_DATA_TEMPR121[17] , \R_DATA_TEMPR121[16] , 
        \R_DATA_TEMPR121[15] , \R_DATA_TEMPR121[14] , 
        \R_DATA_TEMPR121[13] , \R_DATA_TEMPR121[12] , 
        \R_DATA_TEMPR121[11] , \R_DATA_TEMPR121[10] , 
        \R_DATA_TEMPR121[9] , \R_DATA_TEMPR121[8] , 
        \R_DATA_TEMPR121[7] , \R_DATA_TEMPR121[6] , 
        \R_DATA_TEMPR121[5] , \R_DATA_TEMPR121[4] , 
        \R_DATA_TEMPR121[3] , \R_DATA_TEMPR121[2] , 
        \R_DATA_TEMPR121[1] , \R_DATA_TEMPR121[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[121][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[30] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[30] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%18%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C0 (.A_DOUT({
        \R_DATA_TEMPR18[39] , \R_DATA_TEMPR18[38] , 
        \R_DATA_TEMPR18[37] , \R_DATA_TEMPR18[36] , 
        \R_DATA_TEMPR18[35] , \R_DATA_TEMPR18[34] , 
        \R_DATA_TEMPR18[33] , \R_DATA_TEMPR18[32] , 
        \R_DATA_TEMPR18[31] , \R_DATA_TEMPR18[30] , 
        \R_DATA_TEMPR18[29] , \R_DATA_TEMPR18[28] , 
        \R_DATA_TEMPR18[27] , \R_DATA_TEMPR18[26] , 
        \R_DATA_TEMPR18[25] , \R_DATA_TEMPR18[24] , 
        \R_DATA_TEMPR18[23] , \R_DATA_TEMPR18[22] , 
        \R_DATA_TEMPR18[21] , \R_DATA_TEMPR18[20] }), .B_DOUT({
        \R_DATA_TEMPR18[19] , \R_DATA_TEMPR18[18] , 
        \R_DATA_TEMPR18[17] , \R_DATA_TEMPR18[16] , 
        \R_DATA_TEMPR18[15] , \R_DATA_TEMPR18[14] , 
        \R_DATA_TEMPR18[13] , \R_DATA_TEMPR18[12] , 
        \R_DATA_TEMPR18[11] , \R_DATA_TEMPR18[10] , 
        \R_DATA_TEMPR18[9] , \R_DATA_TEMPR18[8] , \R_DATA_TEMPR18[7] , 
        \R_DATA_TEMPR18[6] , \R_DATA_TEMPR18[5] , \R_DATA_TEMPR18[4] , 
        \R_DATA_TEMPR18[3] , \R_DATA_TEMPR18[2] , \R_DATA_TEMPR18[1] , 
        \R_DATA_TEMPR18[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1263 (.A(\R_DATA_TEMPR92[14] ), .B(\R_DATA_TEMPR93[14] ), 
        .C(\R_DATA_TEMPR94[14] ), .D(\R_DATA_TEMPR95[14] ), .Y(
        OR4_1263_Y));
    OR4 OR4_1227 (.A(\R_DATA_TEMPR72[37] ), .B(\R_DATA_TEMPR73[37] ), 
        .C(\R_DATA_TEMPR74[37] ), .D(\R_DATA_TEMPR75[37] ), .Y(
        OR4_1227_Y));
    OR4 OR4_431 (.A(\R_DATA_TEMPR0[7] ), .B(\R_DATA_TEMPR1[7] ), .C(
        \R_DATA_TEMPR2[7] ), .D(\R_DATA_TEMPR3[7] ), .Y(OR4_431_Y));
    OR4 OR4_91 (.A(OR4_893_Y), .B(OR4_692_Y), .C(OR4_349_Y), .D(
        OR4_161_Y), .Y(OR4_91_Y));
    OR4 OR4_1551 (.A(OR4_1291_Y), .B(OR4_1638_Y), .C(OR4_176_Y), .D(
        OR4_1381_Y), .Y(OR4_1551_Y));
    CFG3 #( .INIT(8'h2) )  CFG3_2 (.A(R_EN), .B(R_ADDR[15]), .C(
        R_ADDR[14]), .Y(CFG3_2_Y));
    OR4 OR4_124 (.A(\R_DATA_TEMPR112[31] ), .B(\R_DATA_TEMPR113[31] ), 
        .C(\R_DATA_TEMPR114[31] ), .D(\R_DATA_TEMPR115[31] ), .Y(
        OR4_124_Y));
    OR4 OR4_438 (.A(\R_DATA_TEMPR64[36] ), .B(\R_DATA_TEMPR65[36] ), 
        .C(\R_DATA_TEMPR66[36] ), .D(\R_DATA_TEMPR67[36] ), .Y(
        OR4_438_Y));
    OR4 OR4_1383 (.A(OR4_291_Y), .B(OR4_1591_Y), .C(OR4_1566_Y), .D(
        OR4_925_Y), .Y(OR4_1383_Y));
    OR4 OR4_1030 (.A(OR4_184_Y), .B(OR4_1212_Y), .C(OR4_1473_Y), .D(
        OR4_408_Y), .Y(OR4_1030_Y));
    OR4 OR4_709 (.A(\R_DATA_TEMPR112[24] ), .B(\R_DATA_TEMPR113[24] ), 
        .C(\R_DATA_TEMPR114[24] ), .D(\R_DATA_TEMPR115[24] ), .Y(
        OR4_709_Y));
    OR4 OR4_381 (.A(\R_DATA_TEMPR60[7] ), .B(\R_DATA_TEMPR61[7] ), .C(
        \R_DATA_TEMPR62[7] ), .D(\R_DATA_TEMPR63[7] ), .Y(OR4_381_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[24]  (.A(CFG3_16_Y), .B(
        CFG3_3_Y), .Y(\BLKY2[24] ));
    OR2 OR2_3 (.A(\R_DATA_TEMPR84[13] ), .B(\R_DATA_TEMPR85[13] ), .Y(
        OR2_3_Y));
    OR4 OR4_654 (.A(\R_DATA_TEMPR76[17] ), .B(\R_DATA_TEMPR77[17] ), 
        .C(\R_DATA_TEMPR78[17] ), .D(\R_DATA_TEMPR79[17] ), .Y(
        OR4_654_Y));
    OR4 OR4_947 (.A(\R_DATA_TEMPR80[16] ), .B(\R_DATA_TEMPR81[16] ), 
        .C(\R_DATA_TEMPR82[16] ), .D(\R_DATA_TEMPR83[16] ), .Y(
        OR4_947_Y));
    OR4 OR4_1622 (.A(\R_DATA_TEMPR56[28] ), .B(\R_DATA_TEMPR57[28] ), 
        .C(\R_DATA_TEMPR58[28] ), .D(\R_DATA_TEMPR59[28] ), .Y(
        OR4_1622_Y));
    OR4 OR4_804 (.A(\R_DATA_TEMPR12[25] ), .B(\R_DATA_TEMPR13[25] ), 
        .C(\R_DATA_TEMPR14[25] ), .D(\R_DATA_TEMPR15[25] ), .Y(
        OR4_804_Y));
    OR4 OR4_779 (.A(OR4_83_Y), .B(OR4_1215_Y), .C(OR4_1267_Y), .D(
        OR4_243_Y), .Y(OR4_779_Y));
    OR4 OR4_1426 (.A(\R_DATA_TEMPR80[14] ), .B(\R_DATA_TEMPR81[14] ), 
        .C(\R_DATA_TEMPR82[14] ), .D(\R_DATA_TEMPR83[14] ), .Y(
        OR4_1426_Y));
    OR4 OR4_1324 (.A(\R_DATA_TEMPR120[12] ), .B(\R_DATA_TEMPR121[12] ), 
        .C(\R_DATA_TEMPR122[12] ), .D(\R_DATA_TEMPR123[12] ), .Y(
        OR4_1324_Y));
    OR4 OR4_923 (.A(\R_DATA_TEMPR100[5] ), .B(\R_DATA_TEMPR101[5] ), 
        .C(\R_DATA_TEMPR102[5] ), .D(\R_DATA_TEMPR103[5] ), .Y(
        OR4_923_Y));
    OR4 OR4_480 (.A(\R_DATA_TEMPR40[17] ), .B(\R_DATA_TEMPR41[17] ), 
        .C(\R_DATA_TEMPR42[17] ), .D(\R_DATA_TEMPR43[17] ), .Y(
        OR4_480_Y));
    OR4 OR4_503 (.A(\R_DATA_TEMPR112[20] ), .B(\R_DATA_TEMPR113[20] ), 
        .C(\R_DATA_TEMPR114[20] ), .D(\R_DATA_TEMPR115[20] ), .Y(
        OR4_503_Y));
    OR4 OR4_314 (.A(OR4_1444_Y), .B(OR4_1088_Y), .C(OR4_821_Y), .D(
        OR4_904_Y), .Y(OR4_314_Y));
    CFG3 #( .INIT(8'h80) )  CFG3_21 (.A(R_ADDR[13]), .B(R_ADDR[12]), 
        .C(R_ADDR[11]), .Y(CFG3_21_Y));
    OR4 OR4_1006 (.A(OR4_266_Y), .B(OR4_1432_Y), .C(OR4_341_Y), .D(
        OR4_1360_Y), .Y(OR4_1006_Y));
    OR4 OR4_874 (.A(\R_DATA_TEMPR124[30] ), .B(\R_DATA_TEMPR125[30] ), 
        .C(\R_DATA_TEMPR126[30] ), .D(\R_DATA_TEMPR127[30] ), .Y(
        OR4_874_Y));
    OR4 OR4_826 (.A(\R_DATA_TEMPR100[17] ), .B(\R_DATA_TEMPR101[17] ), 
        .C(\R_DATA_TEMPR102[17] ), .D(\R_DATA_TEMPR103[17] ), .Y(
        OR4_826_Y));
    OR4 OR4_1439 (.A(\R_DATA_TEMPR28[39] ), .B(\R_DATA_TEMPR29[39] ), 
        .C(\R_DATA_TEMPR30[39] ), .D(\R_DATA_TEMPR31[39] ), .Y(
        OR4_1439_Y));
    OR4 OR4_721 (.A(\R_DATA_TEMPR124[31] ), .B(\R_DATA_TEMPR125[31] ), 
        .C(\R_DATA_TEMPR126[31] ), .D(\R_DATA_TEMPR127[31] ), .Y(
        OR4_721_Y));
    OR4 OR4_43 (.A(\R_DATA_TEMPR72[17] ), .B(\R_DATA_TEMPR73[17] ), .C(
        \R_DATA_TEMPR74[17] ), .D(\R_DATA_TEMPR75[17] ), .Y(OR4_43_Y));
    OR4 OR4_1169 (.A(OR4_495_Y), .B(OR4_1056_Y), .C(OR4_1606_Y), .D(
        OR4_425_Y), .Y(OR4_1169_Y));
    OR4 OR4_573 (.A(\R_DATA_TEMPR76[39] ), .B(\R_DATA_TEMPR77[39] ), 
        .C(\R_DATA_TEMPR78[39] ), .D(\R_DATA_TEMPR79[39] ), .Y(
        OR4_573_Y));
    OR4 OR4_539 (.A(\R_DATA_TEMPR16[22] ), .B(\R_DATA_TEMPR17[22] ), 
        .C(\R_DATA_TEMPR18[22] ), .D(\R_DATA_TEMPR19[22] ), .Y(
        OR4_539_Y));
    CFG1 #( .INIT(2'h1) )  \INVBLKX0[0]  (.A(W_ADDR[9]), .Y(\BLKX0[0] )
        );
    OR2 OR2_26 (.A(\R_DATA_TEMPR84[27] ), .B(\R_DATA_TEMPR85[27] ), .Y(
        OR2_26_Y));
    OR4 OR4_111 (.A(\R_DATA_TEMPR32[6] ), .B(\R_DATA_TEMPR33[6] ), .C(
        \R_DATA_TEMPR34[6] ), .D(\R_DATA_TEMPR35[6] ), .Y(OR4_111_Y));
    OR4 OR4_598 (.A(\R_DATA_TEMPR0[25] ), .B(\R_DATA_TEMPR1[25] ), .C(
        \R_DATA_TEMPR2[25] ), .D(\R_DATA_TEMPR3[25] ), .Y(OR4_598_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_1 (.A(R_ADDR[13]), .B(R_ADDR[12]), .C(
        R_ADDR[11]), .Y(CFG3_1_Y));
    OR4 OR4_1627 (.A(\R_DATA_TEMPR100[7] ), .B(\R_DATA_TEMPR101[7] ), 
        .C(\R_DATA_TEMPR102[7] ), .D(\R_DATA_TEMPR103[7] ), .Y(
        OR4_1627_Y));
    OR4 OR4_59 (.A(\R_DATA_TEMPR24[5] ), .B(\R_DATA_TEMPR25[5] ), .C(
        \R_DATA_TEMPR26[5] ), .D(\R_DATA_TEMPR27[5] ), .Y(OR4_59_Y));
    OR4 OR4_530 (.A(\R_DATA_TEMPR116[19] ), .B(\R_DATA_TEMPR117[19] ), 
        .C(\R_DATA_TEMPR118[19] ), .D(\R_DATA_TEMPR119[19] ), .Y(
        OR4_530_Y));
    OR4 OR4_1301 (.A(\R_DATA_TEMPR52[38] ), .B(\R_DATA_TEMPR53[38] ), 
        .C(\R_DATA_TEMPR54[38] ), .D(\R_DATA_TEMPR55[38] ), .Y(
        OR4_1301_Y));
    OR4 OR4_263 (.A(\R_DATA_TEMPR12[26] ), .B(\R_DATA_TEMPR13[26] ), 
        .C(\R_DATA_TEMPR14[26] ), .D(\R_DATA_TEMPR15[26] ), .Y(
        OR4_263_Y));
    OR4 OR4_526 (.A(\R_DATA_TEMPR44[2] ), .B(\R_DATA_TEMPR45[2] ), .C(
        \R_DATA_TEMPR46[2] ), .D(\R_DATA_TEMPR47[2] ), .Y(OR4_526_Y));
    OR4 OR4_1293 (.A(\R_DATA_TEMPR40[3] ), .B(\R_DATA_TEMPR41[3] ), .C(
        \R_DATA_TEMPR42[3] ), .D(\R_DATA_TEMPR43[3] ), .Y(OR4_1293_Y));
    OR4 OR4_1145 (.A(\R_DATA_TEMPR56[5] ), .B(\R_DATA_TEMPR57[5] ), .C(
        \R_DATA_TEMPR58[5] ), .D(\R_DATA_TEMPR59[5] ), .Y(OR4_1145_Y));
    OR4 OR4_445 (.A(OR4_477_Y), .B(OR4_1615_Y), .C(OR4_21_Y), .D(
        OR4_305_Y), .Y(OR4_445_Y));
    OR4 OR4_1329 (.A(OR4_1351_Y), .B(OR4_298_Y), .C(OR4_1072_Y), .D(
        OR4_1338_Y), .Y(OR4_1329_Y));
    OR4 OR4_411 (.A(\R_DATA_TEMPR32[29] ), .B(\R_DATA_TEMPR33[29] ), 
        .C(\R_DATA_TEMPR34[29] ), .D(\R_DATA_TEMPR35[29] ), .Y(
        OR4_411_Y));
    OR4 OR4_1041 (.A(\R_DATA_TEMPR92[10] ), .B(\R_DATA_TEMPR93[10] ), 
        .C(\R_DATA_TEMPR94[10] ), .D(\R_DATA_TEMPR95[10] ), .Y(
        OR4_1041_Y));
    CFG3 #( .INIT(8'h20) )  CFG3_11 (.A(R_ADDR[13]), .B(R_ADDR[12]), 
        .C(R_ADDR[11]), .Y(CFG3_11_Y));
    OR4 OR4_496 (.A(OR4_1424_Y), .B(OR4_238_Y), .C(OR4_1197_Y), .D(
        OR4_1510_Y), .Y(OR4_496_Y));
    OR4 OR4_418 (.A(\R_DATA_TEMPR80[26] ), .B(\R_DATA_TEMPR81[26] ), 
        .C(\R_DATA_TEMPR82[26] ), .D(\R_DATA_TEMPR83[26] ), .Y(
        OR4_418_Y));
    OR4 OR4_1086 (.A(\R_DATA_TEMPR112[7] ), .B(\R_DATA_TEMPR113[7] ), 
        .C(\R_DATA_TEMPR114[7] ), .D(\R_DATA_TEMPR115[7] ), .Y(
        OR4_1086_Y));
    OR4 OR4_1020 (.A(\R_DATA_TEMPR36[27] ), .B(\R_DATA_TEMPR37[27] ), 
        .C(\R_DATA_TEMPR38[27] ), .D(\R_DATA_TEMPR39[27] ), .Y(
        OR4_1020_Y));
    OR4 OR4_968 (.A(\R_DATA_TEMPR108[37] ), .B(\R_DATA_TEMPR109[37] ), 
        .C(\R_DATA_TEMPR110[37] ), .D(\R_DATA_TEMPR111[37] ), .Y(
        OR4_968_Y));
    OR4 OR4_1166 (.A(\R_DATA_TEMPR76[27] ), .B(\R_DATA_TEMPR77[27] ), 
        .C(\R_DATA_TEMPR78[27] ), .D(\R_DATA_TEMPR79[27] ), .Y(
        OR4_1166_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%59%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R59C0 (.A_DOUT({
        \R_DATA_TEMPR59[39] , \R_DATA_TEMPR59[38] , 
        \R_DATA_TEMPR59[37] , \R_DATA_TEMPR59[36] , 
        \R_DATA_TEMPR59[35] , \R_DATA_TEMPR59[34] , 
        \R_DATA_TEMPR59[33] , \R_DATA_TEMPR59[32] , 
        \R_DATA_TEMPR59[31] , \R_DATA_TEMPR59[30] , 
        \R_DATA_TEMPR59[29] , \R_DATA_TEMPR59[28] , 
        \R_DATA_TEMPR59[27] , \R_DATA_TEMPR59[26] , 
        \R_DATA_TEMPR59[25] , \R_DATA_TEMPR59[24] , 
        \R_DATA_TEMPR59[23] , \R_DATA_TEMPR59[22] , 
        \R_DATA_TEMPR59[21] , \R_DATA_TEMPR59[20] }), .B_DOUT({
        \R_DATA_TEMPR59[19] , \R_DATA_TEMPR59[18] , 
        \R_DATA_TEMPR59[17] , \R_DATA_TEMPR59[16] , 
        \R_DATA_TEMPR59[15] , \R_DATA_TEMPR59[14] , 
        \R_DATA_TEMPR59[13] , \R_DATA_TEMPR59[12] , 
        \R_DATA_TEMPR59[11] , \R_DATA_TEMPR59[10] , 
        \R_DATA_TEMPR59[9] , \R_DATA_TEMPR59[8] , \R_DATA_TEMPR59[7] , 
        \R_DATA_TEMPR59[6] , \R_DATA_TEMPR59[5] , \R_DATA_TEMPR59[4] , 
        \R_DATA_TEMPR59[3] , \R_DATA_TEMPR59[2] , \R_DATA_TEMPR59[1] , 
        \R_DATA_TEMPR59[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[59][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[14] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[14] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1461 (.A(\R_DATA_TEMPR88[25] ), .B(\R_DATA_TEMPR89[25] ), 
        .C(\R_DATA_TEMPR90[25] ), .D(\R_DATA_TEMPR91[25] ), .Y(
        OR4_1461_Y));
    OR4 OR4_1381 (.A(OR4_334_Y), .B(OR4_631_Y), .C(OR4_876_Y), .D(
        OR4_678_Y), .Y(OR4_1381_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%62%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R62C0 (.A_DOUT({
        \R_DATA_TEMPR62[39] , \R_DATA_TEMPR62[38] , 
        \R_DATA_TEMPR62[37] , \R_DATA_TEMPR62[36] , 
        \R_DATA_TEMPR62[35] , \R_DATA_TEMPR62[34] , 
        \R_DATA_TEMPR62[33] , \R_DATA_TEMPR62[32] , 
        \R_DATA_TEMPR62[31] , \R_DATA_TEMPR62[30] , 
        \R_DATA_TEMPR62[29] , \R_DATA_TEMPR62[28] , 
        \R_DATA_TEMPR62[27] , \R_DATA_TEMPR62[26] , 
        \R_DATA_TEMPR62[25] , \R_DATA_TEMPR62[24] , 
        \R_DATA_TEMPR62[23] , \R_DATA_TEMPR62[22] , 
        \R_DATA_TEMPR62[21] , \R_DATA_TEMPR62[20] }), .B_DOUT({
        \R_DATA_TEMPR62[19] , \R_DATA_TEMPR62[18] , 
        \R_DATA_TEMPR62[17] , \R_DATA_TEMPR62[16] , 
        \R_DATA_TEMPR62[15] , \R_DATA_TEMPR62[14] , 
        \R_DATA_TEMPR62[13] , \R_DATA_TEMPR62[12] , 
        \R_DATA_TEMPR62[11] , \R_DATA_TEMPR62[10] , 
        \R_DATA_TEMPR62[9] , \R_DATA_TEMPR62[8] , \R_DATA_TEMPR62[7] , 
        \R_DATA_TEMPR62[6] , \R_DATA_TEMPR62[5] , \R_DATA_TEMPR62[4] , 
        \R_DATA_TEMPR62[3] , \R_DATA_TEMPR62[2] , \R_DATA_TEMPR62[1] , 
        \R_DATA_TEMPR62[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[62][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[15] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[15] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[0]  (.A(OR4_1354_Y), .B(OR4_1539_Y), .C(OR4_1016_Y)
        , .D(OR4_1340_Y), .Y(R_DATA[0]));
    OR4 OR4_389 (.A(OR4_929_Y), .B(OR4_1208_Y), .C(OR4_1203_Y), .D(
        OR4_1488_Y), .Y(OR4_389_Y));
    OR4 OR4_1261 (.A(\R_DATA_TEMPR36[24] ), .B(\R_DATA_TEMPR37[24] ), 
        .C(\R_DATA_TEMPR38[24] ), .D(\R_DATA_TEMPR39[24] ), .Y(
        OR4_1261_Y));
    OR4 OR4_392 (.A(\R_DATA_TEMPR52[24] ), .B(\R_DATA_TEMPR53[24] ), 
        .C(\R_DATA_TEMPR54[24] ), .D(\R_DATA_TEMPR55[24] ), .Y(
        OR4_392_Y));
    OR4 OR4_1043 (.A(\R_DATA_TEMPR4[18] ), .B(\R_DATA_TEMPR5[18] ), .C(
        \R_DATA_TEMPR6[18] ), .D(\R_DATA_TEMPR7[18] ), .Y(OR4_1043_Y));
    OR4 OR4_1578 (.A(\R_DATA_TEMPR124[0] ), .B(\R_DATA_TEMPR125[0] ), 
        .C(\R_DATA_TEMPR126[0] ), .D(\R_DATA_TEMPR127[0] ), .Y(
        OR4_1578_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%17%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C0 (.A_DOUT({
        \R_DATA_TEMPR17[39] , \R_DATA_TEMPR17[38] , 
        \R_DATA_TEMPR17[37] , \R_DATA_TEMPR17[36] , 
        \R_DATA_TEMPR17[35] , \R_DATA_TEMPR17[34] , 
        \R_DATA_TEMPR17[33] , \R_DATA_TEMPR17[32] , 
        \R_DATA_TEMPR17[31] , \R_DATA_TEMPR17[30] , 
        \R_DATA_TEMPR17[29] , \R_DATA_TEMPR17[28] , 
        \R_DATA_TEMPR17[27] , \R_DATA_TEMPR17[26] , 
        \R_DATA_TEMPR17[25] , \R_DATA_TEMPR17[24] , 
        \R_DATA_TEMPR17[23] , \R_DATA_TEMPR17[22] , 
        \R_DATA_TEMPR17[21] , \R_DATA_TEMPR17[20] }), .B_DOUT({
        \R_DATA_TEMPR17[19] , \R_DATA_TEMPR17[18] , 
        \R_DATA_TEMPR17[17] , \R_DATA_TEMPR17[16] , 
        \R_DATA_TEMPR17[15] , \R_DATA_TEMPR17[14] , 
        \R_DATA_TEMPR17[13] , \R_DATA_TEMPR17[12] , 
        \R_DATA_TEMPR17[11] , \R_DATA_TEMPR17[10] , 
        \R_DATA_TEMPR17[9] , \R_DATA_TEMPR17[8] , \R_DATA_TEMPR17[7] , 
        \R_DATA_TEMPR17[6] , \R_DATA_TEMPR17[5] , \R_DATA_TEMPR17[4] , 
        \R_DATA_TEMPR17[3] , \R_DATA_TEMPR17[2] , \R_DATA_TEMPR17[1] , 
        \R_DATA_TEMPR17[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%49%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R49C0 (.A_DOUT({
        \R_DATA_TEMPR49[39] , \R_DATA_TEMPR49[38] , 
        \R_DATA_TEMPR49[37] , \R_DATA_TEMPR49[36] , 
        \R_DATA_TEMPR49[35] , \R_DATA_TEMPR49[34] , 
        \R_DATA_TEMPR49[33] , \R_DATA_TEMPR49[32] , 
        \R_DATA_TEMPR49[31] , \R_DATA_TEMPR49[30] , 
        \R_DATA_TEMPR49[29] , \R_DATA_TEMPR49[28] , 
        \R_DATA_TEMPR49[27] , \R_DATA_TEMPR49[26] , 
        \R_DATA_TEMPR49[25] , \R_DATA_TEMPR49[24] , 
        \R_DATA_TEMPR49[23] , \R_DATA_TEMPR49[22] , 
        \R_DATA_TEMPR49[21] , \R_DATA_TEMPR49[20] }), .B_DOUT({
        \R_DATA_TEMPR49[19] , \R_DATA_TEMPR49[18] , 
        \R_DATA_TEMPR49[17] , \R_DATA_TEMPR49[16] , 
        \R_DATA_TEMPR49[15] , \R_DATA_TEMPR49[14] , 
        \R_DATA_TEMPR49[13] , \R_DATA_TEMPR49[12] , 
        \R_DATA_TEMPR49[11] , \R_DATA_TEMPR49[10] , 
        \R_DATA_TEMPR49[9] , \R_DATA_TEMPR49[8] , \R_DATA_TEMPR49[7] , 
        \R_DATA_TEMPR49[6] , \R_DATA_TEMPR49[5] , \R_DATA_TEMPR49[4] , 
        \R_DATA_TEMPR49[3] , \R_DATA_TEMPR49[2] , \R_DATA_TEMPR49[1] , 
        \R_DATA_TEMPR49[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[49][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[12] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[12] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1168 (.A(\R_DATA_TEMPR40[8] ), .B(\R_DATA_TEMPR41[8] ), .C(
        \R_DATA_TEMPR42[8] ), .D(\R_DATA_TEMPR43[8] ), .Y(OR4_1168_Y));
    OR4 OR4_1199 (.A(\R_DATA_TEMPR28[2] ), .B(\R_DATA_TEMPR29[2] ), .C(
        \R_DATA_TEMPR30[2] ), .D(\R_DATA_TEMPR31[2] ), .Y(OR4_1199_Y));
    OR4 OR4_19 (.A(\R_DATA_TEMPR104[38] ), .B(\R_DATA_TEMPR105[38] ), 
        .C(\R_DATA_TEMPR106[38] ), .D(\R_DATA_TEMPR107[38] ), .Y(
        OR4_19_Y));
    OR4 OR4_1429 (.A(OR4_329_Y), .B(OR4_138_Y), .C(OR4_283_Y), .D(
        OR4_1464_Y), .Y(OR4_1429_Y));
    OR4 OR4_41 (.A(\R_DATA_TEMPR64[37] ), .B(\R_DATA_TEMPR65[37] ), .C(
        \R_DATA_TEMPR66[37] ), .D(\R_DATA_TEMPR67[37] ), .Y(OR4_41_Y));
    OR4 OR4_333 (.A(\R_DATA_TEMPR116[25] ), .B(\R_DATA_TEMPR117[25] ), 
        .C(\R_DATA_TEMPR118[25] ), .D(\R_DATA_TEMPR119[25] ), .Y(
        OR4_333_Y));
    OR4 OR4_1442 (.A(\R_DATA_TEMPR60[24] ), .B(\R_DATA_TEMPR61[24] ), 
        .C(\R_DATA_TEMPR62[24] ), .D(\R_DATA_TEMPR63[24] ), .Y(
        OR4_1442_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%38%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R38C0 (.A_DOUT({
        \R_DATA_TEMPR38[39] , \R_DATA_TEMPR38[38] , 
        \R_DATA_TEMPR38[37] , \R_DATA_TEMPR38[36] , 
        \R_DATA_TEMPR38[35] , \R_DATA_TEMPR38[34] , 
        \R_DATA_TEMPR38[33] , \R_DATA_TEMPR38[32] , 
        \R_DATA_TEMPR38[31] , \R_DATA_TEMPR38[30] , 
        \R_DATA_TEMPR38[29] , \R_DATA_TEMPR38[28] , 
        \R_DATA_TEMPR38[27] , \R_DATA_TEMPR38[26] , 
        \R_DATA_TEMPR38[25] , \R_DATA_TEMPR38[24] , 
        \R_DATA_TEMPR38[23] , \R_DATA_TEMPR38[22] , 
        \R_DATA_TEMPR38[21] , \R_DATA_TEMPR38[20] }), .B_DOUT({
        \R_DATA_TEMPR38[19] , \R_DATA_TEMPR38[18] , 
        \R_DATA_TEMPR38[17] , \R_DATA_TEMPR38[16] , 
        \R_DATA_TEMPR38[15] , \R_DATA_TEMPR38[14] , 
        \R_DATA_TEMPR38[13] , \R_DATA_TEMPR38[12] , 
        \R_DATA_TEMPR38[11] , \R_DATA_TEMPR38[10] , 
        \R_DATA_TEMPR38[9] , \R_DATA_TEMPR38[8] , \R_DATA_TEMPR38[7] , 
        \R_DATA_TEMPR38[6] , \R_DATA_TEMPR38[5] , \R_DATA_TEMPR38[4] , 
        \R_DATA_TEMPR38[3] , \R_DATA_TEMPR38[2] , \R_DATA_TEMPR38[1] , 
        \R_DATA_TEMPR38[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[38][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[9] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[9] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_730 (.A(\R_DATA_TEMPR16[28] ), .B(\R_DATA_TEMPR17[28] ), 
        .C(\R_DATA_TEMPR18[28] ), .D(\R_DATA_TEMPR19[28] ), .Y(
        OR4_730_Y));
    OR4 OR4_519 (.A(OR4_1391_Y), .B(OR2_13_Y), .C(\R_DATA_TEMPR86[18] )
        , .D(\R_DATA_TEMPR87[18] ), .Y(OR4_519_Y));
    OR4 OR4_1430 (.A(\R_DATA_TEMPR68[0] ), .B(\R_DATA_TEMPR69[0] ), .C(
        \R_DATA_TEMPR70[0] ), .D(\R_DATA_TEMPR71[0] ), .Y(OR4_1430_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%114%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R114C0 (.A_DOUT({
        \R_DATA_TEMPR114[39] , \R_DATA_TEMPR114[38] , 
        \R_DATA_TEMPR114[37] , \R_DATA_TEMPR114[36] , 
        \R_DATA_TEMPR114[35] , \R_DATA_TEMPR114[34] , 
        \R_DATA_TEMPR114[33] , \R_DATA_TEMPR114[32] , 
        \R_DATA_TEMPR114[31] , \R_DATA_TEMPR114[30] , 
        \R_DATA_TEMPR114[29] , \R_DATA_TEMPR114[28] , 
        \R_DATA_TEMPR114[27] , \R_DATA_TEMPR114[26] , 
        \R_DATA_TEMPR114[25] , \R_DATA_TEMPR114[24] , 
        \R_DATA_TEMPR114[23] , \R_DATA_TEMPR114[22] , 
        \R_DATA_TEMPR114[21] , \R_DATA_TEMPR114[20] }), .B_DOUT({
        \R_DATA_TEMPR114[19] , \R_DATA_TEMPR114[18] , 
        \R_DATA_TEMPR114[17] , \R_DATA_TEMPR114[16] , 
        \R_DATA_TEMPR114[15] , \R_DATA_TEMPR114[14] , 
        \R_DATA_TEMPR114[13] , \R_DATA_TEMPR114[12] , 
        \R_DATA_TEMPR114[11] , \R_DATA_TEMPR114[10] , 
        \R_DATA_TEMPR114[9] , \R_DATA_TEMPR114[8] , 
        \R_DATA_TEMPR114[7] , \R_DATA_TEMPR114[6] , 
        \R_DATA_TEMPR114[5] , \R_DATA_TEMPR114[4] , 
        \R_DATA_TEMPR114[3] , \R_DATA_TEMPR114[2] , 
        \R_DATA_TEMPR114[1] , \R_DATA_TEMPR114[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[114][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[28] , R_ADDR[10], \BLKY0[0] }), 
        .A_CLK(CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], 
        W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], 
        W_DATA[31], W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], 
        W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], 
        W_DATA[21], W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], 
        WBYTE_EN[2]}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], 
        W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], 
        W_ADDR[0], GND, GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[28] , 
        W_ADDR[10], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA[19], 
        W_DATA[18], W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], 
        W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], W_DATA[9], 
        W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], 
        W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1279 (.A(OR4_432_Y), .B(OR4_262_Y), .C(OR4_1285_Y), .D(
        OR4_168_Y), .Y(OR4_1279_Y));
    OR4 OR4_668 (.A(\R_DATA_TEMPR16[33] ), .B(\R_DATA_TEMPR17[33] ), 
        .C(\R_DATA_TEMPR18[33] ), .D(\R_DATA_TEMPR19[33] ), .Y(
        OR4_668_Y));
    OR4 OR4_1613 (.A(\R_DATA_TEMPR96[4] ), .B(\R_DATA_TEMPR97[4] ), .C(
        \R_DATA_TEMPR98[4] ), .D(\R_DATA_TEMPR99[4] ), .Y(OR4_1613_Y));
    OR4 OR4_510 (.A(\R_DATA_TEMPR32[5] ), .B(\R_DATA_TEMPR33[5] ), .C(
        \R_DATA_TEMPR34[5] ), .D(\R_DATA_TEMPR35[5] ), .Y(OR4_510_Y));
    OR4 OR4_1054 (.A(\R_DATA_TEMPR56[9] ), .B(\R_DATA_TEMPR57[9] ), .C(
        \R_DATA_TEMPR58[9] ), .D(\R_DATA_TEMPR59[9] ), .Y(OR4_1054_Y));
    OR4 OR4_432 (.A(\R_DATA_TEMPR96[32] ), .B(\R_DATA_TEMPR97[32] ), 
        .C(\R_DATA_TEMPR98[32] ), .D(\R_DATA_TEMPR99[32] ), .Y(
        OR4_432_Y));
    OR4 OR4_444 (.A(\R_DATA_TEMPR32[7] ), .B(\R_DATA_TEMPR33[7] ), .C(
        \R_DATA_TEMPR34[7] ), .D(\R_DATA_TEMPR35[7] ), .Y(OR4_444_Y));
    OR4 OR4_528 (.A(\R_DATA_TEMPR96[17] ), .B(\R_DATA_TEMPR97[17] ), 
        .C(\R_DATA_TEMPR98[17] ), .D(\R_DATA_TEMPR99[17] ), .Y(
        OR4_528_Y));
    OR4 OR4_52 (.A(\R_DATA_TEMPR68[19] ), .B(\R_DATA_TEMPR69[19] ), .C(
        \R_DATA_TEMPR70[19] ), .D(\R_DATA_TEMPR71[19] ), .Y(OR4_52_Y));
    OR4 OR4_1353 (.A(\R_DATA_TEMPR60[10] ), .B(\R_DATA_TEMPR61[10] ), 
        .C(\R_DATA_TEMPR62[10] ), .D(\R_DATA_TEMPR63[10] ), .Y(
        OR4_1353_Y));
    OR4 OR4_1131 (.A(OR4_306_Y), .B(OR4_1455_Y), .C(OR4_1524_Y), .D(
        OR4_181_Y), .Y(OR4_1131_Y));
    OR4 OR4_662 (.A(\R_DATA_TEMPR32[34] ), .B(\R_DATA_TEMPR33[34] ), 
        .C(\R_DATA_TEMPR34[34] ), .D(\R_DATA_TEMPR35[34] ), .Y(
        OR4_662_Y));
    OR4 OR4_439 (.A(\R_DATA_TEMPR44[7] ), .B(\R_DATA_TEMPR45[7] ), .C(
        \R_DATA_TEMPR46[7] ), .D(\R_DATA_TEMPR47[7] ), .Y(OR4_439_Y));
    OR4 OR4_1514 (.A(OR4_265_Y), .B(OR4_248_Y), .C(OR4_783_Y), .D(
        OR4_177_Y), .Y(OR4_1514_Y));
    CFG3 #( .INIT(8'h2) )  CFG3_18 (.A(R_ADDR[13]), .B(R_ADDR[12]), .C(
        R_ADDR[11]), .Y(CFG3_18_Y));
    OR4 OR4_346 (.A(\R_DATA_TEMPR20[38] ), .B(\R_DATA_TEMPR21[38] ), 
        .C(\R_DATA_TEMPR22[38] ), .D(\R_DATA_TEMPR23[38] ), .Y(
        OR4_346_Y));
    OR2 OR2_20 (.A(\R_DATA_TEMPR84[0] ), .B(\R_DATA_TEMPR85[0] ), .Y(
        OR2_20_Y));
    OR4 OR4_136 (.A(\R_DATA_TEMPR116[39] ), .B(\R_DATA_TEMPR117[39] ), 
        .C(\R_DATA_TEMPR118[39] ), .D(\R_DATA_TEMPR119[39] ), .Y(
        OR4_136_Y));
    CFG1 #( .INIT(2'h1) )  \INVBLKX1[0]  (.A(W_ADDR[10]), .Y(
        \BLKX1[0] ));
    OR4 OR4_1315 (.A(OR4_1607_Y), .B(OR4_551_Y), .C(OR4_1337_Y), .D(
        OR4_1597_Y), .Y(OR4_1315_Y));
    OR4 OR4_1536 (.A(\R_DATA_TEMPR56[23] ), .B(\R_DATA_TEMPR57[23] ), 
        .C(\R_DATA_TEMPR58[23] ), .D(\R_DATA_TEMPR59[23] ), .Y(
        OR4_1536_Y));
    OR2 OR2_16 (.A(\R_DATA_TEMPR84[32] ), .B(\R_DATA_TEMPR85[32] ), .Y(
        OR2_16_Y));
    CFG3 #( .INIT(8'h20) )  CFG3_22 (.A(W_ADDR[13]), .B(W_ADDR[12]), 
        .C(W_ADDR[11]), .Y(CFG3_22_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[20]  (.A(CFG3_18_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[20] ));
    OR2 OR2_27 (.A(\R_DATA_TEMPR84[19] ), .B(\R_DATA_TEMPR85[19] ), .Y(
        OR2_27_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%55%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R55C0 (.A_DOUT({
        \R_DATA_TEMPR55[39] , \R_DATA_TEMPR55[38] , 
        \R_DATA_TEMPR55[37] , \R_DATA_TEMPR55[36] , 
        \R_DATA_TEMPR55[35] , \R_DATA_TEMPR55[34] , 
        \R_DATA_TEMPR55[33] , \R_DATA_TEMPR55[32] , 
        \R_DATA_TEMPR55[31] , \R_DATA_TEMPR55[30] , 
        \R_DATA_TEMPR55[29] , \R_DATA_TEMPR55[28] , 
        \R_DATA_TEMPR55[27] , \R_DATA_TEMPR55[26] , 
        \R_DATA_TEMPR55[25] , \R_DATA_TEMPR55[24] , 
        \R_DATA_TEMPR55[23] , \R_DATA_TEMPR55[22] , 
        \R_DATA_TEMPR55[21] , \R_DATA_TEMPR55[20] }), .B_DOUT({
        \R_DATA_TEMPR55[19] , \R_DATA_TEMPR55[18] , 
        \R_DATA_TEMPR55[17] , \R_DATA_TEMPR55[16] , 
        \R_DATA_TEMPR55[15] , \R_DATA_TEMPR55[14] , 
        \R_DATA_TEMPR55[13] , \R_DATA_TEMPR55[12] , 
        \R_DATA_TEMPR55[11] , \R_DATA_TEMPR55[10] , 
        \R_DATA_TEMPR55[9] , \R_DATA_TEMPR55[8] , \R_DATA_TEMPR55[7] , 
        \R_DATA_TEMPR55[6] , \R_DATA_TEMPR55[5] , \R_DATA_TEMPR55[4] , 
        \R_DATA_TEMPR55[3] , \R_DATA_TEMPR55[2] , \R_DATA_TEMPR55[1] , 
        \R_DATA_TEMPR55[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[55][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[13] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[13] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_426 (.A(OR4_169_Y), .B(OR4_750_Y), .C(OR4_1536_Y), .D(
        OR4_155_Y), .Y(OR4_426_Y));
    OR4 OR4_1196 (.A(OR4_1602_Y), .B(OR4_278_Y), .C(OR4_524_Y), .D(
        OR4_337_Y), .Y(OR4_1196_Y));
    OR4 OR4_203 (.A(OR4_901_Y), .B(OR4_569_Y), .C(OR4_1090_Y), .D(
        OR4_1545_Y), .Y(OR4_203_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[19]  (.A(CFG3_5_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[19] ));
    OR4 OR4_290 (.A(\R_DATA_TEMPR100[4] ), .B(\R_DATA_TEMPR101[4] ), 
        .C(\R_DATA_TEMPR102[4] ), .D(\R_DATA_TEMPR103[4] ), .Y(
        OR4_290_Y));
    OR4 OR4_1491 (.A(OR4_69_Y), .B(OR4_850_Y), .C(OR4_1319_Y), .D(
        OR4_1626_Y), .Y(OR4_1491_Y));
    OR4 OR4_597 (.A(OR4_101_Y), .B(OR4_412_Y), .C(OR4_650_Y), .D(
        OR4_464_Y), .Y(OR4_597_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%45%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R45C0 (.A_DOUT({
        \R_DATA_TEMPR45[39] , \R_DATA_TEMPR45[38] , 
        \R_DATA_TEMPR45[37] , \R_DATA_TEMPR45[36] , 
        \R_DATA_TEMPR45[35] , \R_DATA_TEMPR45[34] , 
        \R_DATA_TEMPR45[33] , \R_DATA_TEMPR45[32] , 
        \R_DATA_TEMPR45[31] , \R_DATA_TEMPR45[30] , 
        \R_DATA_TEMPR45[29] , \R_DATA_TEMPR45[28] , 
        \R_DATA_TEMPR45[27] , \R_DATA_TEMPR45[26] , 
        \R_DATA_TEMPR45[25] , \R_DATA_TEMPR45[24] , 
        \R_DATA_TEMPR45[23] , \R_DATA_TEMPR45[22] , 
        \R_DATA_TEMPR45[21] , \R_DATA_TEMPR45[20] }), .B_DOUT({
        \R_DATA_TEMPR45[19] , \R_DATA_TEMPR45[18] , 
        \R_DATA_TEMPR45[17] , \R_DATA_TEMPR45[16] , 
        \R_DATA_TEMPR45[15] , \R_DATA_TEMPR45[14] , 
        \R_DATA_TEMPR45[13] , \R_DATA_TEMPR45[12] , 
        \R_DATA_TEMPR45[11] , \R_DATA_TEMPR45[10] , 
        \R_DATA_TEMPR45[9] , \R_DATA_TEMPR45[8] , \R_DATA_TEMPR45[7] , 
        \R_DATA_TEMPR45[6] , \R_DATA_TEMPR45[5] , \R_DATA_TEMPR45[4] , 
        \R_DATA_TEMPR45[3] , \R_DATA_TEMPR45[2] , \R_DATA_TEMPR45[1] , 
        \R_DATA_TEMPR45[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[45][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[11] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[11] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1102 (.A(\R_DATA_TEMPR20[15] ), .B(\R_DATA_TEMPR21[15] ), 
        .C(\R_DATA_TEMPR22[15] ), .D(\R_DATA_TEMPR23[15] ), .Y(
        OR4_1102_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%92%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R92C0 (.A_DOUT({
        \R_DATA_TEMPR92[39] , \R_DATA_TEMPR92[38] , 
        \R_DATA_TEMPR92[37] , \R_DATA_TEMPR92[36] , 
        \R_DATA_TEMPR92[35] , \R_DATA_TEMPR92[34] , 
        \R_DATA_TEMPR92[33] , \R_DATA_TEMPR92[32] , 
        \R_DATA_TEMPR92[31] , \R_DATA_TEMPR92[30] , 
        \R_DATA_TEMPR92[29] , \R_DATA_TEMPR92[28] , 
        \R_DATA_TEMPR92[27] , \R_DATA_TEMPR92[26] , 
        \R_DATA_TEMPR92[25] , \R_DATA_TEMPR92[24] , 
        \R_DATA_TEMPR92[23] , \R_DATA_TEMPR92[22] , 
        \R_DATA_TEMPR92[21] , \R_DATA_TEMPR92[20] }), .B_DOUT({
        \R_DATA_TEMPR92[19] , \R_DATA_TEMPR92[18] , 
        \R_DATA_TEMPR92[17] , \R_DATA_TEMPR92[16] , 
        \R_DATA_TEMPR92[15] , \R_DATA_TEMPR92[14] , 
        \R_DATA_TEMPR92[13] , \R_DATA_TEMPR92[12] , 
        \R_DATA_TEMPR92[11] , \R_DATA_TEMPR92[10] , 
        \R_DATA_TEMPR92[9] , \R_DATA_TEMPR92[8] , \R_DATA_TEMPR92[7] , 
        \R_DATA_TEMPR92[6] , \R_DATA_TEMPR92[5] , \R_DATA_TEMPR92[4] , 
        \R_DATA_TEMPR92[3] , \R_DATA_TEMPR92[2] , \R_DATA_TEMPR92[1] , 
        \R_DATA_TEMPR92[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[92][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[23] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[23] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1291 (.A(OR4_1540_Y), .B(OR4_686_Y), .C(OR4_1144_Y), .D(
        OR4_1481_Y), .Y(OR4_1291_Y));
    OR4 OR4_858 (.A(OR4_146_Y), .B(OR2_15_Y), .C(\R_DATA_TEMPR86[8] ), 
        .D(\R_DATA_TEMPR87[8] ), .Y(OR4_858_Y));
    OR4 OR4_789 (.A(\R_DATA_TEMPR88[9] ), .B(\R_DATA_TEMPR89[9] ), .C(
        \R_DATA_TEMPR90[9] ), .D(\R_DATA_TEMPR91[9] ), .Y(OR4_789_Y));
    OR4 OR4_338 (.A(OR4_191_Y), .B(OR4_456_Y), .C(OR4_635_Y), .D(
        OR4_340_Y), .Y(OR4_338_Y));
    OR4 OR4_273 (.A(\R_DATA_TEMPR0[18] ), .B(\R_DATA_TEMPR1[18] ), .C(
        \R_DATA_TEMPR2[18] ), .D(\R_DATA_TEMPR3[18] ), .Y(OR4_273_Y));
    OR4 OR4_1198 (.A(OR4_354_Y), .B(OR4_1026_Y), .C(OR4_1580_Y), .D(
        OR4_970_Y), .Y(OR4_1198_Y));
    OR4 OR4_908 (.A(OR4_1092_Y), .B(OR4_977_Y), .C(OR4_1518_Y), .D(
        OR4_351_Y), .Y(OR4_908_Y));
    OR4 OR4_1437 (.A(\R_DATA_TEMPR80[29] ), .B(\R_DATA_TEMPR81[29] ), 
        .C(\R_DATA_TEMPR82[29] ), .D(\R_DATA_TEMPR83[29] ), .Y(
        OR4_1437_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%113%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R113C0 (.A_DOUT({
        \R_DATA_TEMPR113[39] , \R_DATA_TEMPR113[38] , 
        \R_DATA_TEMPR113[37] , \R_DATA_TEMPR113[36] , 
        \R_DATA_TEMPR113[35] , \R_DATA_TEMPR113[34] , 
        \R_DATA_TEMPR113[33] , \R_DATA_TEMPR113[32] , 
        \R_DATA_TEMPR113[31] , \R_DATA_TEMPR113[30] , 
        \R_DATA_TEMPR113[29] , \R_DATA_TEMPR113[28] , 
        \R_DATA_TEMPR113[27] , \R_DATA_TEMPR113[26] , 
        \R_DATA_TEMPR113[25] , \R_DATA_TEMPR113[24] , 
        \R_DATA_TEMPR113[23] , \R_DATA_TEMPR113[22] , 
        \R_DATA_TEMPR113[21] , \R_DATA_TEMPR113[20] }), .B_DOUT({
        \R_DATA_TEMPR113[19] , \R_DATA_TEMPR113[18] , 
        \R_DATA_TEMPR113[17] , \R_DATA_TEMPR113[16] , 
        \R_DATA_TEMPR113[15] , \R_DATA_TEMPR113[14] , 
        \R_DATA_TEMPR113[13] , \R_DATA_TEMPR113[12] , 
        \R_DATA_TEMPR113[11] , \R_DATA_TEMPR113[10] , 
        \R_DATA_TEMPR113[9] , \R_DATA_TEMPR113[8] , 
        \R_DATA_TEMPR113[7] , \R_DATA_TEMPR113[6] , 
        \R_DATA_TEMPR113[5] , \R_DATA_TEMPR113[4] , 
        \R_DATA_TEMPR113[3] , \R_DATA_TEMPR113[2] , 
        \R_DATA_TEMPR113[1] , \R_DATA_TEMPR113[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[113][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[28] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[28] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_313 (.A(\R_DATA_TEMPR36[20] ), .B(\R_DATA_TEMPR37[20] ), 
        .C(\R_DATA_TEMPR38[20] ), .D(\R_DATA_TEMPR39[20] ), .Y(
        OR4_313_Y));
    OR4 OR4_322 (.A(OR4_68_Y), .B(OR4_1447_Y), .C(OR4_1137_Y), .D(
        OR4_1290_Y), .Y(OR4_322_Y));
    OR4 OR4_865 (.A(OR4_1416_Y), .B(OR4_1069_Y), .C(OR4_1045_Y), .D(
        OR4_426_Y), .Y(OR4_865_Y));
    OR4 OR4_710 (.A(\R_DATA_TEMPR100[31] ), .B(\R_DATA_TEMPR101[31] ), 
        .C(\R_DATA_TEMPR102[31] ), .D(\R_DATA_TEMPR103[31] ), .Y(
        OR4_710_Y));
    OR4 OR4_1420 (.A(\R_DATA_TEMPR68[34] ), .B(\R_DATA_TEMPR69[34] ), 
        .C(\R_DATA_TEMPR70[34] ), .D(\R_DATA_TEMPR71[34] ), .Y(
        OR4_1420_Y));
    OR4 OR4_1048 (.A(\R_DATA_TEMPR12[15] ), .B(\R_DATA_TEMPR13[15] ), 
        .C(\R_DATA_TEMPR14[15] ), .D(\R_DATA_TEMPR15[15] ), .Y(
        OR4_1048_Y));
    OR4 OR4_884 (.A(\R_DATA_TEMPR124[3] ), .B(\R_DATA_TEMPR125[3] ), 
        .C(\R_DATA_TEMPR126[3] ), .D(\R_DATA_TEMPR127[3] ), .Y(
        OR4_884_Y));
    OR4 OR4_699 (.A(\R_DATA_TEMPR0[31] ), .B(\R_DATA_TEMPR1[31] ), .C(
        \R_DATA_TEMPR2[31] ), .D(\R_DATA_TEMPR3[31] ), .Y(OR4_699_Y));
    OR4 OR4_12 (.A(\R_DATA_TEMPR28[16] ), .B(\R_DATA_TEMPR29[16] ), .C(
        \R_DATA_TEMPR30[16] ), .D(\R_DATA_TEMPR31[16] ), .Y(OR4_12_Y));
    OR4 OR4_978 (.A(\R_DATA_TEMPR12[4] ), .B(\R_DATA_TEMPR13[4] ), .C(
        \R_DATA_TEMPR14[4] ), .D(\R_DATA_TEMPR15[4] ), .Y(OR4_978_Y));
    CFG3 #( .INIT(8'h2) )  CFG3_12 (.A(W_EN), .B(W_ADDR[15]), .C(
        W_ADDR[14]), .Y(CFG3_12_Y));
    OR4 OR4_583 (.A(\R_DATA_TEMPR104[22] ), .B(\R_DATA_TEMPR105[22] ), 
        .C(\R_DATA_TEMPR106[22] ), .D(\R_DATA_TEMPR107[22] ), .Y(
        OR4_583_Y));
    OR4 OR4_412 (.A(\R_DATA_TEMPR100[18] ), .B(\R_DATA_TEMPR101[18] ), 
        .C(\R_DATA_TEMPR102[18] ), .D(\R_DATA_TEMPR103[18] ), .Y(
        OR4_412_Y));
    OR4 OR4_1035 (.A(\R_DATA_TEMPR124[8] ), .B(\R_DATA_TEMPR125[8] ), 
        .C(\R_DATA_TEMPR126[8] ), .D(\R_DATA_TEMPR127[8] ), .Y(
        OR4_1035_Y));
    OR4 OR4_296 (.A(\R_DATA_TEMPR80[5] ), .B(\R_DATA_TEMPR81[5] ), .C(
        \R_DATA_TEMPR82[5] ), .D(\R_DATA_TEMPR83[5] ), .Y(OR4_296_Y));
    OR4 OR4_1121 (.A(\R_DATA_TEMPR124[26] ), .B(\R_DATA_TEMPR125[26] ), 
        .C(\R_DATA_TEMPR126[26] ), .D(\R_DATA_TEMPR127[26] ), .Y(
        OR4_1121_Y));
    OR4 OR4_1056 (.A(\R_DATA_TEMPR36[0] ), .B(\R_DATA_TEMPR37[0] ), .C(
        \R_DATA_TEMPR38[0] ), .D(\R_DATA_TEMPR39[0] ), .Y(OR4_1056_Y));
    OR4 OR4_419 (.A(\R_DATA_TEMPR108[35] ), .B(\R_DATA_TEMPR109[35] ), 
        .C(\R_DATA_TEMPR110[35] ), .D(\R_DATA_TEMPR111[35] ), .Y(
        OR4_419_Y));
    OR4 OR4_251 (.A(OR4_1151_Y), .B(OR4_1430_Y), .C(OR4_1611_Y), .D(
        OR4_1382_Y), .Y(OR4_251_Y));
    OR4 OR4_79 (.A(\R_DATA_TEMPR52[7] ), .B(\R_DATA_TEMPR53[7] ), .C(
        \R_DATA_TEMPR54[7] ), .D(\R_DATA_TEMPR55[7] ), .Y(OR4_79_Y));
    OR4 OR4_1542 (.A(\R_DATA_TEMPR104[29] ), .B(\R_DATA_TEMPR105[29] ), 
        .C(\R_DATA_TEMPR106[29] ), .D(\R_DATA_TEMPR107[29] ), .Y(
        OR4_1542_Y));
    CFG3 #( .INIT(8'h40) )  CFG3_19 (.A(R_ADDR[13]), .B(R_ADDR[12]), 
        .C(R_ADDR[11]), .Y(CFG3_19_Y));
    OR4 OR4_139 (.A(\R_DATA_TEMPR56[39] ), .B(\R_DATA_TEMPR57[39] ), 
        .C(\R_DATA_TEMPR58[39] ), .D(\R_DATA_TEMPR59[39] ), .Y(
        OR4_139_Y));
    OR4 OR4_116 (.A(\R_DATA_TEMPR64[11] ), .B(\R_DATA_TEMPR65[11] ), 
        .C(\R_DATA_TEMPR66[11] ), .D(\R_DATA_TEMPR67[11] ), .Y(
        OR4_116_Y));
    OR4 OR4_1182 (.A(\R_DATA_TEMPR108[9] ), .B(\R_DATA_TEMPR109[9] ), 
        .C(\R_DATA_TEMPR110[9] ), .D(\R_DATA_TEMPR111[9] ), .Y(
        OR4_1182_Y));
    OR4 OR4_608 (.A(OR4_1162_Y), .B(OR4_1492_Y), .C(OR4_928_Y), .D(
        OR4_141_Y), .Y(OR4_608_Y));
    OR4 OR4_144 (.A(\R_DATA_TEMPR112[23] ), .B(\R_DATA_TEMPR113[23] ), 
        .C(\R_DATA_TEMPR114[23] ), .D(\R_DATA_TEMPR115[23] ), .Y(
        OR4_144_Y));
    OR4 OR4_1526 (.A(\R_DATA_TEMPR124[7] ), .B(\R_DATA_TEMPR125[7] ), 
        .C(\R_DATA_TEMPR126[7] ), .D(\R_DATA_TEMPR127[7] ), .Y(
        OR4_1526_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%37%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R37C0 (.A_DOUT({
        \R_DATA_TEMPR37[39] , \R_DATA_TEMPR37[38] , 
        \R_DATA_TEMPR37[37] , \R_DATA_TEMPR37[36] , 
        \R_DATA_TEMPR37[35] , \R_DATA_TEMPR37[34] , 
        \R_DATA_TEMPR37[33] , \R_DATA_TEMPR37[32] , 
        \R_DATA_TEMPR37[31] , \R_DATA_TEMPR37[30] , 
        \R_DATA_TEMPR37[29] , \R_DATA_TEMPR37[28] , 
        \R_DATA_TEMPR37[27] , \R_DATA_TEMPR37[26] , 
        \R_DATA_TEMPR37[25] , \R_DATA_TEMPR37[24] , 
        \R_DATA_TEMPR37[23] , \R_DATA_TEMPR37[22] , 
        \R_DATA_TEMPR37[21] , \R_DATA_TEMPR37[20] }), .B_DOUT({
        \R_DATA_TEMPR37[19] , \R_DATA_TEMPR37[18] , 
        \R_DATA_TEMPR37[17] , \R_DATA_TEMPR37[16] , 
        \R_DATA_TEMPR37[15] , \R_DATA_TEMPR37[14] , 
        \R_DATA_TEMPR37[13] , \R_DATA_TEMPR37[12] , 
        \R_DATA_TEMPR37[11] , \R_DATA_TEMPR37[10] , 
        \R_DATA_TEMPR37[9] , \R_DATA_TEMPR37[8] , \R_DATA_TEMPR37[7] , 
        \R_DATA_TEMPR37[6] , \R_DATA_TEMPR37[5] , \R_DATA_TEMPR37[4] , 
        \R_DATA_TEMPR37[3] , \R_DATA_TEMPR37[2] , \R_DATA_TEMPR37[1] , 
        \R_DATA_TEMPR37[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[37][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[9] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[9] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_694 (.A(\R_DATA_TEMPR24[35] ), .B(\R_DATA_TEMPR25[35] ), 
        .C(\R_DATA_TEMPR26[35] ), .D(\R_DATA_TEMPR27[35] ), .Y(
        OR4_694_Y));
    OR4 OR4_1351 (.A(\R_DATA_TEMPR48[29] ), .B(\R_DATA_TEMPR49[29] ), 
        .C(\R_DATA_TEMPR50[29] ), .D(\R_DATA_TEMPR51[29] ), .Y(
        OR4_1351_Y));
    OR4 OR4_678 (.A(\R_DATA_TEMPR60[14] ), .B(\R_DATA_TEMPR61[14] ), 
        .C(\R_DATA_TEMPR62[14] ), .D(\R_DATA_TEMPR63[14] ), .Y(
        OR4_678_Y));
    OR4 OR4_602 (.A(OR4_0_Y), .B(OR2_22_Y), .C(\R_DATA_TEMPR86[11] ), 
        .D(\R_DATA_TEMPR87[11] ), .Y(OR4_602_Y));
    OR4 \OR4_R_DATA[32]  (.A(OR4_1557_Y), .B(OR4_1512_Y), .C(
        OR4_1279_Y), .D(OR4_556_Y), .Y(R_DATA[32]));
    OR4 OR4_552 (.A(\R_DATA_TEMPR28[26] ), .B(\R_DATA_TEMPR29[26] ), 
        .C(\R_DATA_TEMPR30[26] ), .D(\R_DATA_TEMPR31[26] ), .Y(
        OR4_552_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[25]  (.A(CFG3_8_Y), .B(CFG3_7_Y)
        , .Y(\BLKX2[25] ));
    OR4 OR4_931 (.A(OR4_623_Y), .B(OR2_34_Y), .C(\R_DATA_TEMPR86[17] ), 
        .D(\R_DATA_TEMPR87[17] ), .Y(OR4_931_Y));
    OR4 OR4_943 (.A(\R_DATA_TEMPR24[2] ), .B(\R_DATA_TEMPR25[2] ), .C(
        \R_DATA_TEMPR26[2] ), .D(\R_DATA_TEMPR27[2] ), .Y(OR4_943_Y));
    OR4 OR4_220 (.A(\R_DATA_TEMPR80[31] ), .B(\R_DATA_TEMPR81[31] ), 
        .C(\R_DATA_TEMPR82[31] ), .D(\R_DATA_TEMPR83[31] ), .Y(
        OR4_220_Y));
    OR4 OR4_1273 (.A(\R_DATA_TEMPR12[35] ), .B(\R_DATA_TEMPR13[35] ), 
        .C(\R_DATA_TEMPR14[35] ), .D(\R_DATA_TEMPR15[35] ), .Y(
        OR4_1273_Y));
    OR4 OR4_672 (.A(\R_DATA_TEMPR68[24] ), .B(\R_DATA_TEMPR69[24] ), 
        .C(\R_DATA_TEMPR70[24] ), .D(\R_DATA_TEMPR71[24] ), .Y(
        OR4_672_Y));
    OR4 OR4_527 (.A(OR4_1167_Y), .B(OR4_91_Y), .C(OR4_787_Y), .D(
        OR4_1471_Y), .Y(OR4_527_Y));
    OR4 OR4_318 (.A(\R_DATA_TEMPR28[0] ), .B(\R_DATA_TEMPR29[0] ), .C(
        \R_DATA_TEMPR30[0] ), .D(\R_DATA_TEMPR31[0] ), .Y(OR4_318_Y));
    OR2 OR2_10 (.A(\R_DATA_TEMPR84[15] ), .B(\R_DATA_TEMPR85[15] ), .Y(
        OR2_10_Y));
    OR4 OR4_846 (.A(\R_DATA_TEMPR120[5] ), .B(\R_DATA_TEMPR121[5] ), 
        .C(\R_DATA_TEMPR122[5] ), .D(\R_DATA_TEMPR123[5] ), .Y(
        OR4_846_Y));
    OR4 OR4_1427 (.A(\R_DATA_TEMPR4[10] ), .B(\R_DATA_TEMPR5[10] ), .C(
        \R_DATA_TEMPR6[10] ), .D(\R_DATA_TEMPR7[10] ), .Y(OR4_1427_Y));
    OR4 OR4_741 (.A(OR4_500_Y), .B(OR4_942_Y), .C(OR4_288_Y), .D(
        OR4_592_Y), .Y(OR4_741_Y));
    OR4 OR4_1012 (.A(OR4_1209_Y), .B(OR4_142_Y), .C(OR4_934_Y), .D(
        OR4_1192_Y), .Y(OR4_1012_Y));
    OR4 \OR4_R_DATA[3]  (.A(OR4_398_Y), .B(OR4_847_Y), .C(OR4_718_Y), 
        .D(OR4_843_Y), .Y(R_DATA[3]));
    OR2 OR2_17 (.A(\R_DATA_TEMPR84[2] ), .B(\R_DATA_TEMPR85[2] ), .Y(
        OR2_17_Y));
    OR4 OR4_666 (.A(\R_DATA_TEMPR96[35] ), .B(\R_DATA_TEMPR97[35] ), 
        .C(\R_DATA_TEMPR98[35] ), .D(\R_DATA_TEMPR99[35] ), .Y(
        OR4_666_Y));
    OR4 OR4_629 (.A(\R_DATA_TEMPR12[31] ), .B(\R_DATA_TEMPR13[31] ), 
        .C(\R_DATA_TEMPR14[31] ), .D(\R_DATA_TEMPR15[31] ), .Y(
        OR4_629_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%76%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R76C0 (.A_DOUT({
        \R_DATA_TEMPR76[39] , \R_DATA_TEMPR76[38] , 
        \R_DATA_TEMPR76[37] , \R_DATA_TEMPR76[36] , 
        \R_DATA_TEMPR76[35] , \R_DATA_TEMPR76[34] , 
        \R_DATA_TEMPR76[33] , \R_DATA_TEMPR76[32] , 
        \R_DATA_TEMPR76[31] , \R_DATA_TEMPR76[30] , 
        \R_DATA_TEMPR76[29] , \R_DATA_TEMPR76[28] , 
        \R_DATA_TEMPR76[27] , \R_DATA_TEMPR76[26] , 
        \R_DATA_TEMPR76[25] , \R_DATA_TEMPR76[24] , 
        \R_DATA_TEMPR76[23] , \R_DATA_TEMPR76[22] , 
        \R_DATA_TEMPR76[21] , \R_DATA_TEMPR76[20] }), .B_DOUT({
        \R_DATA_TEMPR76[19] , \R_DATA_TEMPR76[18] , 
        \R_DATA_TEMPR76[17] , \R_DATA_TEMPR76[16] , 
        \R_DATA_TEMPR76[15] , \R_DATA_TEMPR76[14] , 
        \R_DATA_TEMPR76[13] , \R_DATA_TEMPR76[12] , 
        \R_DATA_TEMPR76[11] , \R_DATA_TEMPR76[10] , 
        \R_DATA_TEMPR76[9] , \R_DATA_TEMPR76[8] , \R_DATA_TEMPR76[7] , 
        \R_DATA_TEMPR76[6] , \R_DATA_TEMPR76[5] , \R_DATA_TEMPR76[4] , 
        \R_DATA_TEMPR76[3] , \R_DATA_TEMPR76[2] , \R_DATA_TEMPR76[1] , 
        \R_DATA_TEMPR76[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[76][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[19] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[19] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1025 (.A(OR4_882_Y), .B(OR2_9_Y), .C(\R_DATA_TEMPR86[24] ), 
        .D(\R_DATA_TEMPR87[24] ), .Y(OR4_1025_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%110%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R110C0 (.A_DOUT({
        \R_DATA_TEMPR110[39] , \R_DATA_TEMPR110[38] , 
        \R_DATA_TEMPR110[37] , \R_DATA_TEMPR110[36] , 
        \R_DATA_TEMPR110[35] , \R_DATA_TEMPR110[34] , 
        \R_DATA_TEMPR110[33] , \R_DATA_TEMPR110[32] , 
        \R_DATA_TEMPR110[31] , \R_DATA_TEMPR110[30] , 
        \R_DATA_TEMPR110[29] , \R_DATA_TEMPR110[28] , 
        \R_DATA_TEMPR110[27] , \R_DATA_TEMPR110[26] , 
        \R_DATA_TEMPR110[25] , \R_DATA_TEMPR110[24] , 
        \R_DATA_TEMPR110[23] , \R_DATA_TEMPR110[22] , 
        \R_DATA_TEMPR110[21] , \R_DATA_TEMPR110[20] }), .B_DOUT({
        \R_DATA_TEMPR110[19] , \R_DATA_TEMPR110[18] , 
        \R_DATA_TEMPR110[17] , \R_DATA_TEMPR110[16] , 
        \R_DATA_TEMPR110[15] , \R_DATA_TEMPR110[14] , 
        \R_DATA_TEMPR110[13] , \R_DATA_TEMPR110[12] , 
        \R_DATA_TEMPR110[11] , \R_DATA_TEMPR110[10] , 
        \R_DATA_TEMPR110[9] , \R_DATA_TEMPR110[8] , 
        \R_DATA_TEMPR110[7] , \R_DATA_TEMPR110[6] , 
        \R_DATA_TEMPR110[5] , \R_DATA_TEMPR110[4] , 
        \R_DATA_TEMPR110[3] , \R_DATA_TEMPR110[2] , 
        \R_DATA_TEMPR110[1] , \R_DATA_TEMPR110[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[110][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[27] , R_ADDR[10], \BLKY0[0] }), 
        .A_CLK(CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], 
        W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], 
        W_DATA[31], W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], 
        W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], 
        W_DATA[21], W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], 
        WBYTE_EN[2]}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], 
        W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], 
        W_ADDR[0], GND, GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[27] , 
        W_ADDR[10], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA[19], 
        W_DATA[18], W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], 
        W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], W_DATA[9], 
        W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], 
        W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%19%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C0 (.A_DOUT({
        \R_DATA_TEMPR19[39] , \R_DATA_TEMPR19[38] , 
        \R_DATA_TEMPR19[37] , \R_DATA_TEMPR19[36] , 
        \R_DATA_TEMPR19[35] , \R_DATA_TEMPR19[34] , 
        \R_DATA_TEMPR19[33] , \R_DATA_TEMPR19[32] , 
        \R_DATA_TEMPR19[31] , \R_DATA_TEMPR19[30] , 
        \R_DATA_TEMPR19[29] , \R_DATA_TEMPR19[28] , 
        \R_DATA_TEMPR19[27] , \R_DATA_TEMPR19[26] , 
        \R_DATA_TEMPR19[25] , \R_DATA_TEMPR19[24] , 
        \R_DATA_TEMPR19[23] , \R_DATA_TEMPR19[22] , 
        \R_DATA_TEMPR19[21] , \R_DATA_TEMPR19[20] }), .B_DOUT({
        \R_DATA_TEMPR19[19] , \R_DATA_TEMPR19[18] , 
        \R_DATA_TEMPR19[17] , \R_DATA_TEMPR19[16] , 
        \R_DATA_TEMPR19[15] , \R_DATA_TEMPR19[14] , 
        \R_DATA_TEMPR19[13] , \R_DATA_TEMPR19[12] , 
        \R_DATA_TEMPR19[11] , \R_DATA_TEMPR19[10] , 
        \R_DATA_TEMPR19[9] , \R_DATA_TEMPR19[8] , \R_DATA_TEMPR19[7] , 
        \R_DATA_TEMPR19[6] , \R_DATA_TEMPR19[5] , \R_DATA_TEMPR19[4] , 
        \R_DATA_TEMPR19[3] , \R_DATA_TEMPR19[2] , \R_DATA_TEMPR19[1] , 
        \R_DATA_TEMPR19[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_554 (.A(\R_DATA_TEMPR108[38] ), .B(\R_DATA_TEMPR109[38] ), 
        .C(\R_DATA_TEMPR110[38] ), .D(\R_DATA_TEMPR111[38] ), .Y(
        OR4_554_Y));
    OR4 OR4_952 (.A(\R_DATA_TEMPR8[30] ), .B(\R_DATA_TEMPR9[30] ), .C(
        \R_DATA_TEMPR10[30] ), .D(\R_DATA_TEMPR11[30] ), .Y(OR4_952_Y));
    OR4 OR4_546 (.A(\R_DATA_TEMPR88[29] ), .B(\R_DATA_TEMPR89[29] ), 
        .C(\R_DATA_TEMPR90[29] ), .D(\R_DATA_TEMPR91[29] ), .Y(
        OR4_546_Y));
    OR4 OR4_226 (.A(\R_DATA_TEMPR76[25] ), .B(\R_DATA_TEMPR77[25] ), 
        .C(\R_DATA_TEMPR78[25] ), .D(\R_DATA_TEMPR79[25] ), .Y(
        OR4_226_Y));
    OR4 OR4_119 (.A(\R_DATA_TEMPR0[34] ), .B(\R_DATA_TEMPR1[34] ), .C(
        \R_DATA_TEMPR2[34] ), .D(\R_DATA_TEMPR3[34] ), .Y(OR4_119_Y));
    OR4 OR4_1047 (.A(\R_DATA_TEMPR116[35] ), .B(\R_DATA_TEMPR117[35] ), 
        .C(\R_DATA_TEMPR118[35] ), .D(\R_DATA_TEMPR119[35] ), .Y(
        OR4_1047_Y));
    OR4 OR4_805 (.A(\R_DATA_TEMPR12[23] ), .B(\R_DATA_TEMPR13[23] ), 
        .C(\R_DATA_TEMPR14[23] ), .D(\R_DATA_TEMPR15[23] ), .Y(
        OR4_805_Y));
    OR4 OR4_1179 (.A(\R_DATA_TEMPR48[36] ), .B(\R_DATA_TEMPR49[36] ), 
        .C(\R_DATA_TEMPR50[36] ), .D(\R_DATA_TEMPR51[36] ), .Y(
        OR4_1179_Y));
    OR4 OR4_72 (.A(\R_DATA_TEMPR100[33] ), .B(\R_DATA_TEMPR101[33] ), 
        .C(\R_DATA_TEMPR102[33] ), .D(\R_DATA_TEMPR103[33] ), .Y(
        OR4_72_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%86%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R86C0 (.A_DOUT({
        \R_DATA_TEMPR86[39] , \R_DATA_TEMPR86[38] , 
        \R_DATA_TEMPR86[37] , \R_DATA_TEMPR86[36] , 
        \R_DATA_TEMPR86[35] , \R_DATA_TEMPR86[34] , 
        \R_DATA_TEMPR86[33] , \R_DATA_TEMPR86[32] , 
        \R_DATA_TEMPR86[31] , \R_DATA_TEMPR86[30] , 
        \R_DATA_TEMPR86[29] , \R_DATA_TEMPR86[28] , 
        \R_DATA_TEMPR86[27] , \R_DATA_TEMPR86[26] , 
        \R_DATA_TEMPR86[25] , \R_DATA_TEMPR86[24] , 
        \R_DATA_TEMPR86[23] , \R_DATA_TEMPR86[22] , 
        \R_DATA_TEMPR86[21] , \R_DATA_TEMPR86[20] }), .B_DOUT({
        \R_DATA_TEMPR86[19] , \R_DATA_TEMPR86[18] , 
        \R_DATA_TEMPR86[17] , \R_DATA_TEMPR86[16] , 
        \R_DATA_TEMPR86[15] , \R_DATA_TEMPR86[14] , 
        \R_DATA_TEMPR86[13] , \R_DATA_TEMPR86[12] , 
        \R_DATA_TEMPR86[11] , \R_DATA_TEMPR86[10] , 
        \R_DATA_TEMPR86[9] , \R_DATA_TEMPR86[8] , \R_DATA_TEMPR86[7] , 
        \R_DATA_TEMPR86[6] , \R_DATA_TEMPR86[5] , \R_DATA_TEMPR86[4] , 
        \R_DATA_TEMPR86[3] , \R_DATA_TEMPR86[2] , \R_DATA_TEMPR86[1] , 
        \R_DATA_TEMPR86[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[86][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[21] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[21] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1130 (.A(\R_DATA_TEMPR28[12] ), .B(\R_DATA_TEMPR29[12] ), 
        .C(\R_DATA_TEMPR30[12] ), .D(\R_DATA_TEMPR31[12] ), .Y(
        OR4_1130_Y));
    OR4 OR4_875 (.A(OR4_218_Y), .B(OR4_52_Y), .C(OR4_175_Y), .D(
        OR4_369_Y), .Y(OR4_875_Y));
    OR4 OR4_735 (.A(\R_DATA_TEMPR36[14] ), .B(\R_DATA_TEMPR37[14] ), 
        .C(\R_DATA_TEMPR38[14] ), .D(\R_DATA_TEMPR39[14] ), .Y(
        OR4_735_Y));
    OR4 OR4_637 (.A(\R_DATA_TEMPR56[4] ), .B(\R_DATA_TEMPR57[4] ), .C(
        \R_DATA_TEMPR58[4] ), .D(\R_DATA_TEMPR59[4] ), .Y(OR4_637_Y));
    OR4 OR4_736 (.A(\R_DATA_TEMPR24[13] ), .B(\R_DATA_TEMPR25[13] ), 
        .C(\R_DATA_TEMPR26[13] ), .D(\R_DATA_TEMPR27[13] ), .Y(
        OR4_736_Y));
    OR4 OR4_624 (.A(\R_DATA_TEMPR100[34] ), .B(\R_DATA_TEMPR101[34] ), 
        .C(\R_DATA_TEMPR102[34] ), .D(\R_DATA_TEMPR103[34] ), .Y(
        OR4_624_Y));
    OR4 OR4_1564 (.A(\R_DATA_TEMPR44[23] ), .B(\R_DATA_TEMPR45[23] ), 
        .C(\R_DATA_TEMPR46[23] ), .D(\R_DATA_TEMPR47[23] ), .Y(
        OR4_1564_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[30]  (.A(CFG3_10_Y), .B(
        CFG3_7_Y), .Y(\BLKX2[30] ));
    OR4 OR4_351 (.A(\R_DATA_TEMPR44[9] ), .B(\R_DATA_TEMPR45[9] ), .C(
        \R_DATA_TEMPR46[9] ), .D(\R_DATA_TEMPR47[9] ), .Y(OR4_351_Y));
    OR2 OR2_28 (.A(\R_DATA_TEMPR84[35] ), .B(\R_DATA_TEMPR85[35] ), .Y(
        OR2_28_Y));
    OR4 \OR4_R_DATA[33]  (.A(OR4_1383_Y), .B(OR4_941_Y), .C(OR4_890_Y), 
        .D(OR4_827_Y), .Y(R_DATA[33]));
    OR4 OR4_911 (.A(\R_DATA_TEMPR28[9] ), .B(\R_DATA_TEMPR29[9] ), .C(
        \R_DATA_TEMPR30[9] ), .D(\R_DATA_TEMPR31[9] ), .Y(OR4_911_Y));
    OR4 OR4_1365 (.A(OR4_1445_Y), .B(OR2_8_Y), .C(\R_DATA_TEMPR86[1] ), 
        .D(\R_DATA_TEMPR87[1] ), .Y(OR4_1365_Y));
    OR4 OR4_1508 (.A(\R_DATA_TEMPR24[18] ), .B(\R_DATA_TEMPR25[18] ), 
        .C(\R_DATA_TEMPR26[18] ), .D(\R_DATA_TEMPR27[18] ), .Y(
        OR4_1508_Y));
    OR4 \OR4_R_DATA[25]  (.A(OR4_1288_Y), .B(OR4_440_Y), .C(OR4_1059_Y)
        , .D(OR4_605_Y), .Y(R_DATA[25]));
    OR4 OR4_450 (.A(\R_DATA_TEMPR68[30] ), .B(\R_DATA_TEMPR69[30] ), 
        .C(\R_DATA_TEMPR70[30] ), .D(\R_DATA_TEMPR71[30] ), .Y(
        OR4_450_Y));
    OR4 OR4_283 (.A(\R_DATA_TEMPR72[14] ), .B(\R_DATA_TEMPR73[14] ), 
        .C(\R_DATA_TEMPR74[14] ), .D(\R_DATA_TEMPR75[14] ), .Y(
        OR4_283_Y));
    OR4 OR4_96 (.A(\R_DATA_TEMPR104[13] ), .B(\R_DATA_TEMPR105[13] ), 
        .C(\R_DATA_TEMPR106[13] ), .D(\R_DATA_TEMPR107[13] ), .Y(
        OR4_96_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%15%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C0 (.A_DOUT({
        \R_DATA_TEMPR15[39] , \R_DATA_TEMPR15[38] , 
        \R_DATA_TEMPR15[37] , \R_DATA_TEMPR15[36] , 
        \R_DATA_TEMPR15[35] , \R_DATA_TEMPR15[34] , 
        \R_DATA_TEMPR15[33] , \R_DATA_TEMPR15[32] , 
        \R_DATA_TEMPR15[31] , \R_DATA_TEMPR15[30] , 
        \R_DATA_TEMPR15[29] , \R_DATA_TEMPR15[28] , 
        \R_DATA_TEMPR15[27] , \R_DATA_TEMPR15[26] , 
        \R_DATA_TEMPR15[25] , \R_DATA_TEMPR15[24] , 
        \R_DATA_TEMPR15[23] , \R_DATA_TEMPR15[22] , 
        \R_DATA_TEMPR15[21] , \R_DATA_TEMPR15[20] }), .B_DOUT({
        \R_DATA_TEMPR15[19] , \R_DATA_TEMPR15[18] , 
        \R_DATA_TEMPR15[17] , \R_DATA_TEMPR15[16] , 
        \R_DATA_TEMPR15[15] , \R_DATA_TEMPR15[14] , 
        \R_DATA_TEMPR15[13] , \R_DATA_TEMPR15[12] , 
        \R_DATA_TEMPR15[11] , \R_DATA_TEMPR15[10] , 
        \R_DATA_TEMPR15[9] , \R_DATA_TEMPR15[8] , \R_DATA_TEMPR15[7] , 
        \R_DATA_TEMPR15[6] , \R_DATA_TEMPR15[5] , \R_DATA_TEMPR15[4] , 
        \R_DATA_TEMPR15[3] , \R_DATA_TEMPR15[2] , \R_DATA_TEMPR15[1] , 
        \R_DATA_TEMPR15[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1209 (.A(\R_DATA_TEMPR48[27] ), .B(\R_DATA_TEMPR49[27] ), 
        .C(\R_DATA_TEMPR50[27] ), .D(\R_DATA_TEMPR51[27] ), .Y(
        OR4_1209_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_17 (.A(W_EN), .B(W_ADDR[15]), .C(
        W_ADDR[14]), .Y(CFG3_17_Y));
    OR4 OR4_1513 (.A(\R_DATA_TEMPR8[18] ), .B(\R_DATA_TEMPR9[18] ), .C(
        \R_DATA_TEMPR10[18] ), .D(\R_DATA_TEMPR11[18] ), .Y(OR4_1513_Y)
        );
    OR4 OR4_1330 (.A(\R_DATA_TEMPR120[31] ), .B(\R_DATA_TEMPR121[31] ), 
        .C(\R_DATA_TEMPR122[31] ), .D(\R_DATA_TEMPR123[31] ), .Y(
        OR4_1330_Y));
    OR4 OR4_1176 (.A(OR4_1240_Y), .B(OR4_121_Y), .C(OR4_1262_Y), .D(
        OR4_771_Y), .Y(OR4_1176_Y));
    OR4 OR4_548 (.A(\R_DATA_TEMPR36[11] ), .B(\R_DATA_TEMPR37[11] ), 
        .C(\R_DATA_TEMPR38[11] ), .D(\R_DATA_TEMPR39[11] ), .Y(
        OR4_548_Y));
    OR4 OR4_1471 (.A(OR4_227_Y), .B(OR4_541_Y), .C(OR4_776_Y), .D(
        OR4_588_Y), .Y(OR4_1471_Y));
    OR4 OR4_1152 (.A(\R_DATA_TEMPR36[2] ), .B(\R_DATA_TEMPR37[2] ), .C(
        \R_DATA_TEMPR38[2] ), .D(\R_DATA_TEMPR39[2] ), .Y(OR4_1152_Y));
    OR4 OR4_54 (.A(\R_DATA_TEMPR24[31] ), .B(\R_DATA_TEMPR25[31] ), .C(
        \R_DATA_TEMPR26[31] ), .D(\R_DATA_TEMPR27[31] ), .Y(OR4_54_Y));
    OR4 OR4_988 (.A(OR4_767_Y), .B(OR4_1474_Y), .C(OR4_373_Y), .D(
        OR4_1409_Y), .Y(OR4_988_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%112%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R112C0 (.A_DOUT({
        \R_DATA_TEMPR112[39] , \R_DATA_TEMPR112[38] , 
        \R_DATA_TEMPR112[37] , \R_DATA_TEMPR112[36] , 
        \R_DATA_TEMPR112[35] , \R_DATA_TEMPR112[34] , 
        \R_DATA_TEMPR112[33] , \R_DATA_TEMPR112[32] , 
        \R_DATA_TEMPR112[31] , \R_DATA_TEMPR112[30] , 
        \R_DATA_TEMPR112[29] , \R_DATA_TEMPR112[28] , 
        \R_DATA_TEMPR112[27] , \R_DATA_TEMPR112[26] , 
        \R_DATA_TEMPR112[25] , \R_DATA_TEMPR112[24] , 
        \R_DATA_TEMPR112[23] , \R_DATA_TEMPR112[22] , 
        \R_DATA_TEMPR112[21] , \R_DATA_TEMPR112[20] }), .B_DOUT({
        \R_DATA_TEMPR112[19] , \R_DATA_TEMPR112[18] , 
        \R_DATA_TEMPR112[17] , \R_DATA_TEMPR112[16] , 
        \R_DATA_TEMPR112[15] , \R_DATA_TEMPR112[14] , 
        \R_DATA_TEMPR112[13] , \R_DATA_TEMPR112[12] , 
        \R_DATA_TEMPR112[11] , \R_DATA_TEMPR112[10] , 
        \R_DATA_TEMPR112[9] , \R_DATA_TEMPR112[8] , 
        \R_DATA_TEMPR112[7] , \R_DATA_TEMPR112[6] , 
        \R_DATA_TEMPR112[5] , \R_DATA_TEMPR112[4] , 
        \R_DATA_TEMPR112[3] , \R_DATA_TEMPR112[2] , 
        \R_DATA_TEMPR112[1] , \R_DATA_TEMPR112[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[112][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[28] , \BLKY1[0] , \BLKY0[0] }), 
        .A_CLK(CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], 
        W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], 
        W_DATA[31], W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], 
        W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], 
        W_DATA[21], W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], 
        WBYTE_EN[2]}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], 
        W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], 
        W_ADDR[0], GND, GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[28] , 
        \BLKX1[0] , \BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA[19], 
        W_DATA[18], W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], 
        W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], W_DATA[9], 
        W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], 
        W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1271 (.A(\R_DATA_TEMPR52[8] ), .B(\R_DATA_TEMPR53[8] ), .C(
        \R_DATA_TEMPR54[8] ), .D(\R_DATA_TEMPR55[8] ), .Y(OR4_1271_Y));
    OR4 OR4_3 (.A(\R_DATA_TEMPR116[4] ), .B(\R_DATA_TEMPR117[4] ), .C(
        \R_DATA_TEMPR118[4] ), .D(\R_DATA_TEMPR119[4] ), .Y(OR4_3_Y));
    OR4 OR4_1178 (.A(\R_DATA_TEMPR116[38] ), .B(\R_DATA_TEMPR117[38] ), 
        .C(\R_DATA_TEMPR118[38] ), .D(\R_DATA_TEMPR119[38] ), .Y(
        OR4_1178_Y));
    OR4 OR4_364 (.A(\R_DATA_TEMPR88[15] ), .B(\R_DATA_TEMPR89[15] ), 
        .C(\R_DATA_TEMPR90[15] ), .D(\R_DATA_TEMPR91[15] ), .Y(
        OR4_364_Y));
    OR4 OR4_1120 (.A(\R_DATA_TEMPR120[13] ), .B(\R_DATA_TEMPR121[13] ), 
        .C(\R_DATA_TEMPR122[13] ), .D(\R_DATA_TEMPR123[13] ), .Y(
        OR4_1120_Y));
    OR4 OR4_606 (.A(\R_DATA_TEMPR28[20] ), .B(\R_DATA_TEMPR29[20] ), 
        .C(\R_DATA_TEMPR30[20] ), .D(\R_DATA_TEMPR31[20] ), .Y(
        OR4_606_Y));
    OR4 OR4_1588 (.A(OR4_1186_Y), .B(OR4_1465_Y), .C(OR4_951_Y), .D(
        OR4_687_Y), .Y(OR4_1588_Y));
    OR4 OR4_715 (.A(OR4_435_Y), .B(OR4_241_Y), .C(OR4_1508_Y), .D(
        OR4_1346_Y), .Y(OR4_715_Y));
    OR4 OR4_617 (.A(\R_DATA_TEMPR124[22] ), .B(\R_DATA_TEMPR125[22] ), 
        .C(\R_DATA_TEMPR126[22] ), .D(\R_DATA_TEMPR127[22] ), .Y(
        OR4_617_Y));
    OR4 OR4_161 (.A(\R_DATA_TEMPR28[19] ), .B(\R_DATA_TEMPR29[19] ), 
        .C(\R_DATA_TEMPR30[19] ), .D(\R_DATA_TEMPR31[19] ), .Y(
        OR4_161_Y));
    OR4 OR4_446 (.A(OR4_1066_Y), .B(OR4_910_Y), .C(OR4_1023_Y), .D(
        OR4_768_Y), .Y(OR4_446_Y));
    OR4 OR4_1594 (.A(OR4_1007_Y), .B(OR2_3_Y), .C(\R_DATA_TEMPR86[13] )
        , .D(\R_DATA_TEMPR87[13] ), .Y(OR4_1594_Y));
    OR4 OR4_716 (.A(\R_DATA_TEMPR64[38] ), .B(\R_DATA_TEMPR65[38] ), 
        .C(\R_DATA_TEMPR66[38] ), .D(\R_DATA_TEMPR67[38] ), .Y(
        OR4_716_Y));
    OR4 OR4_676 (.A(OR4_7_Y), .B(OR4_1484_Y), .C(OR4_872_Y), .D(
        OR4_1402_Y), .Y(OR4_676_Y));
    OR4 OR4_1289 (.A(\R_DATA_TEMPR92[5] ), .B(\R_DATA_TEMPR93[5] ), .C(
        \R_DATA_TEMPR94[5] ), .D(\R_DATA_TEMPR95[5] ), .Y(OR4_1289_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[6]  (.A(CFG3_1_Y), .B(CFG3_2_Y), 
        .Y(\BLKY2[6] ));
    OR4 OR4_237 (.A(\R_DATA_TEMPR116[20] ), .B(\R_DATA_TEMPR117[20] ), 
        .C(\R_DATA_TEMPR118[20] ), .D(\R_DATA_TEMPR119[20] ), .Y(
        OR4_237_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%39%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R39C0 (.A_DOUT({
        \R_DATA_TEMPR39[39] , \R_DATA_TEMPR39[38] , 
        \R_DATA_TEMPR39[37] , \R_DATA_TEMPR39[36] , 
        \R_DATA_TEMPR39[35] , \R_DATA_TEMPR39[34] , 
        \R_DATA_TEMPR39[33] , \R_DATA_TEMPR39[32] , 
        \R_DATA_TEMPR39[31] , \R_DATA_TEMPR39[30] , 
        \R_DATA_TEMPR39[29] , \R_DATA_TEMPR39[28] , 
        \R_DATA_TEMPR39[27] , \R_DATA_TEMPR39[26] , 
        \R_DATA_TEMPR39[25] , \R_DATA_TEMPR39[24] , 
        \R_DATA_TEMPR39[23] , \R_DATA_TEMPR39[22] , 
        \R_DATA_TEMPR39[21] , \R_DATA_TEMPR39[20] }), .B_DOUT({
        \R_DATA_TEMPR39[19] , \R_DATA_TEMPR39[18] , 
        \R_DATA_TEMPR39[17] , \R_DATA_TEMPR39[16] , 
        \R_DATA_TEMPR39[15] , \R_DATA_TEMPR39[14] , 
        \R_DATA_TEMPR39[13] , \R_DATA_TEMPR39[12] , 
        \R_DATA_TEMPR39[11] , \R_DATA_TEMPR39[10] , 
        \R_DATA_TEMPR39[9] , \R_DATA_TEMPR39[8] , \R_DATA_TEMPR39[7] , 
        \R_DATA_TEMPR39[6] , \R_DATA_TEMPR39[5] , \R_DATA_TEMPR39[4] , 
        \R_DATA_TEMPR39[3] , \R_DATA_TEMPR39[2] , \R_DATA_TEMPR39[1] , 
        \R_DATA_TEMPR39[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[39][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[9] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[9] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_898 (.A(OR4_1063_Y), .B(OR4_506_Y), .C(OR4_1071_Y), .D(
        OR4_455_Y), .Y(OR4_898_Y));
    OR4 OR4_688 (.A(\R_DATA_TEMPR56[38] ), .B(\R_DATA_TEMPR57[38] ), 
        .C(\R_DATA_TEMPR58[38] ), .D(\R_DATA_TEMPR59[38] ), .Y(
        OR4_688_Y));
    OR4 OR4_1395 (.A(\R_DATA_TEMPR112[4] ), .B(\R_DATA_TEMPR113[4] ), 
        .C(\R_DATA_TEMPR114[4] ), .D(\R_DATA_TEMPR115[4] ), .Y(
        OR4_1395_Y));
    OR4 OR4_137 (.A(\R_DATA_TEMPR20[2] ), .B(\R_DATA_TEMPR21[2] ), .C(
        \R_DATA_TEMPR22[2] ), .D(\R_DATA_TEMPR23[2] ), .Y(OR4_137_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%126%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R126C0 (.A_DOUT({
        \R_DATA_TEMPR126[39] , \R_DATA_TEMPR126[38] , 
        \R_DATA_TEMPR126[37] , \R_DATA_TEMPR126[36] , 
        \R_DATA_TEMPR126[35] , \R_DATA_TEMPR126[34] , 
        \R_DATA_TEMPR126[33] , \R_DATA_TEMPR126[32] , 
        \R_DATA_TEMPR126[31] , \R_DATA_TEMPR126[30] , 
        \R_DATA_TEMPR126[29] , \R_DATA_TEMPR126[28] , 
        \R_DATA_TEMPR126[27] , \R_DATA_TEMPR126[26] , 
        \R_DATA_TEMPR126[25] , \R_DATA_TEMPR126[24] , 
        \R_DATA_TEMPR126[23] , \R_DATA_TEMPR126[22] , 
        \R_DATA_TEMPR126[21] , \R_DATA_TEMPR126[20] }), .B_DOUT({
        \R_DATA_TEMPR126[19] , \R_DATA_TEMPR126[18] , 
        \R_DATA_TEMPR126[17] , \R_DATA_TEMPR126[16] , 
        \R_DATA_TEMPR126[15] , \R_DATA_TEMPR126[14] , 
        \R_DATA_TEMPR126[13] , \R_DATA_TEMPR126[12] , 
        \R_DATA_TEMPR126[11] , \R_DATA_TEMPR126[10] , 
        \R_DATA_TEMPR126[9] , \R_DATA_TEMPR126[8] , 
        \R_DATA_TEMPR126[7] , \R_DATA_TEMPR126[6] , 
        \R_DATA_TEMPR126[5] , \R_DATA_TEMPR126[4] , 
        \R_DATA_TEMPR126[3] , \R_DATA_TEMPR126[2] , 
        \R_DATA_TEMPR126[1] , \R_DATA_TEMPR126[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[126][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[31] , R_ADDR[10], \BLKY0[0] }), 
        .A_CLK(CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], 
        W_DATA[36], W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], 
        W_DATA[31], W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], 
        W_DATA[26], W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], 
        W_DATA[21], W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], 
        WBYTE_EN[2]}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], 
        W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], 
        W_ADDR[0], GND, GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[31] , 
        W_ADDR[10], \BLKX0[0] }), .B_CLK(CLK), .B_DIN({W_DATA[19], 
        W_DATA[18], W_DATA[17], W_DATA[16], W_DATA[15], W_DATA[14], 
        W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], W_DATA[9], 
        W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], W_DATA[4], 
        W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), .B_REN(VCC), 
        .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%51%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R51C0 (.A_DOUT({
        \R_DATA_TEMPR51[39] , \R_DATA_TEMPR51[38] , 
        \R_DATA_TEMPR51[37] , \R_DATA_TEMPR51[36] , 
        \R_DATA_TEMPR51[35] , \R_DATA_TEMPR51[34] , 
        \R_DATA_TEMPR51[33] , \R_DATA_TEMPR51[32] , 
        \R_DATA_TEMPR51[31] , \R_DATA_TEMPR51[30] , 
        \R_DATA_TEMPR51[29] , \R_DATA_TEMPR51[28] , 
        \R_DATA_TEMPR51[27] , \R_DATA_TEMPR51[26] , 
        \R_DATA_TEMPR51[25] , \R_DATA_TEMPR51[24] , 
        \R_DATA_TEMPR51[23] , \R_DATA_TEMPR51[22] , 
        \R_DATA_TEMPR51[21] , \R_DATA_TEMPR51[20] }), .B_DOUT({
        \R_DATA_TEMPR51[19] , \R_DATA_TEMPR51[18] , 
        \R_DATA_TEMPR51[17] , \R_DATA_TEMPR51[16] , 
        \R_DATA_TEMPR51[15] , \R_DATA_TEMPR51[14] , 
        \R_DATA_TEMPR51[13] , \R_DATA_TEMPR51[12] , 
        \R_DATA_TEMPR51[11] , \R_DATA_TEMPR51[10] , 
        \R_DATA_TEMPR51[9] , \R_DATA_TEMPR51[8] , \R_DATA_TEMPR51[7] , 
        \R_DATA_TEMPR51[6] , \R_DATA_TEMPR51[5] , \R_DATA_TEMPR51[4] , 
        \R_DATA_TEMPR51[3] , \R_DATA_TEMPR51[2] , \R_DATA_TEMPR51[1] , 
        \R_DATA_TEMPR51[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[51][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[12] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[12] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1235 (.A(OR4_173_Y), .B(OR4_696_Y), .C(OR4_208_Y), .D(
        OR4_1341_Y), .Y(OR4_1235_Y));
    OR4 OR4_682 (.A(\R_DATA_TEMPR108[0] ), .B(\R_DATA_TEMPR109[0] ), 
        .C(\R_DATA_TEMPR110[0] ), .D(\R_DATA_TEMPR111[0] ), .Y(
        OR4_682_Y));
    OR4 OR4_342 (.A(OR4_892_Y), .B(OR4_710_Y), .C(OR4_112_Y), .D(
        OR4_630_Y), .Y(OR4_342_Y));
    OR4 OR4_359 (.A(OR4_944_Y), .B(OR2_16_Y), .C(\R_DATA_TEMPR86[32] ), 
        .D(\R_DATA_TEMPR87[32] ), .Y(OR4_359_Y));
    OR4 OR4_461 (.A(\R_DATA_TEMPR108[14] ), .B(\R_DATA_TEMPR109[14] ), 
        .C(\R_DATA_TEMPR110[14] ), .D(\R_DATA_TEMPR111[14] ), .Y(
        OR4_461_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[11]  (.A(CFG3_5_Y), .B(CFG3_4_Y)
        , .Y(\BLKX2[11] ));
    OR4 OR4_14 (.A(\R_DATA_TEMPR76[34] ), .B(\R_DATA_TEMPR77[34] ), .C(
        \R_DATA_TEMPR78[34] ), .D(\R_DATA_TEMPR79[34] ), .Y(OR4_14_Y));
    OR4 OR4_1531 (.A(\R_DATA_TEMPR108[13] ), .B(\R_DATA_TEMPR109[13] ), 
        .C(\R_DATA_TEMPR110[13] ), .D(\R_DATA_TEMPR111[13] ), .Y(
        OR4_1531_Y));
    OR4 OR4_468 (.A(\R_DATA_TEMPR92[31] ), .B(\R_DATA_TEMPR93[31] ), 
        .C(\R_DATA_TEMPR94[31] ), .D(\R_DATA_TEMPR95[31] ), .Y(
        OR4_468_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%41%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R41C0 (.A_DOUT({
        \R_DATA_TEMPR41[39] , \R_DATA_TEMPR41[38] , 
        \R_DATA_TEMPR41[37] , \R_DATA_TEMPR41[36] , 
        \R_DATA_TEMPR41[35] , \R_DATA_TEMPR41[34] , 
        \R_DATA_TEMPR41[33] , \R_DATA_TEMPR41[32] , 
        \R_DATA_TEMPR41[31] , \R_DATA_TEMPR41[30] , 
        \R_DATA_TEMPR41[29] , \R_DATA_TEMPR41[28] , 
        \R_DATA_TEMPR41[27] , \R_DATA_TEMPR41[26] , 
        \R_DATA_TEMPR41[25] , \R_DATA_TEMPR41[24] , 
        \R_DATA_TEMPR41[23] , \R_DATA_TEMPR41[22] , 
        \R_DATA_TEMPR41[21] , \R_DATA_TEMPR41[20] }), .B_DOUT({
        \R_DATA_TEMPR41[19] , \R_DATA_TEMPR41[18] , 
        \R_DATA_TEMPR41[17] , \R_DATA_TEMPR41[16] , 
        \R_DATA_TEMPR41[15] , \R_DATA_TEMPR41[14] , 
        \R_DATA_TEMPR41[13] , \R_DATA_TEMPR41[12] , 
        \R_DATA_TEMPR41[11] , \R_DATA_TEMPR41[10] , 
        \R_DATA_TEMPR41[9] , \R_DATA_TEMPR41[8] , \R_DATA_TEMPR41[7] , 
        \R_DATA_TEMPR41[6] , \R_DATA_TEMPR41[5] , \R_DATA_TEMPR41[4] , 
        \R_DATA_TEMPR41[3] , \R_DATA_TEMPR41[2] , \R_DATA_TEMPR41[1] , 
        \R_DATA_TEMPR41[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[41][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[10] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[10] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1320 (.A(\R_DATA_TEMPR112[32] ), .B(\R_DATA_TEMPR113[32] ), 
        .C(\R_DATA_TEMPR114[32] ), .D(\R_DATA_TEMPR115[32] ), .Y(
        OR4_1320_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%24%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C0 (.A_DOUT({
        \R_DATA_TEMPR24[39] , \R_DATA_TEMPR24[38] , 
        \R_DATA_TEMPR24[37] , \R_DATA_TEMPR24[36] , 
        \R_DATA_TEMPR24[35] , \R_DATA_TEMPR24[34] , 
        \R_DATA_TEMPR24[33] , \R_DATA_TEMPR24[32] , 
        \R_DATA_TEMPR24[31] , \R_DATA_TEMPR24[30] , 
        \R_DATA_TEMPR24[29] , \R_DATA_TEMPR24[28] , 
        \R_DATA_TEMPR24[27] , \R_DATA_TEMPR24[26] , 
        \R_DATA_TEMPR24[25] , \R_DATA_TEMPR24[24] , 
        \R_DATA_TEMPR24[23] , \R_DATA_TEMPR24[22] , 
        \R_DATA_TEMPR24[21] , \R_DATA_TEMPR24[20] }), .B_DOUT({
        \R_DATA_TEMPR24[19] , \R_DATA_TEMPR24[18] , 
        \R_DATA_TEMPR24[17] , \R_DATA_TEMPR24[16] , 
        \R_DATA_TEMPR24[15] , \R_DATA_TEMPR24[14] , 
        \R_DATA_TEMPR24[13] , \R_DATA_TEMPR24[12] , 
        \R_DATA_TEMPR24[11] , \R_DATA_TEMPR24[10] , 
        \R_DATA_TEMPR24[9] , \R_DATA_TEMPR24[8] , \R_DATA_TEMPR24[7] , 
        \R_DATA_TEMPR24[6] , \R_DATA_TEMPR24[5] , \R_DATA_TEMPR24[4] , 
        \R_DATA_TEMPR24[3] , \R_DATA_TEMPR24[2] , \R_DATA_TEMPR24[1] , 
        \R_DATA_TEMPR24[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR2 OR2_18 (.A(\R_DATA_TEMPR84[30] ), .B(\R_DATA_TEMPR85[30] ), .Y(
        OR2_18_Y));
    OR4 OR4_1247 (.A(\R_DATA_TEMPR104[19] ), .B(\R_DATA_TEMPR105[19] ), 
        .C(\R_DATA_TEMPR106[19] ), .D(\R_DATA_TEMPR107[19] ), .Y(
        OR4_1247_Y));
    OR4 OR4_733 (.A(OR4_844_Y), .B(OR4_585_Y), .C(OR4_303_Y), .D(
        OR4_889_Y), .Y(OR4_733_Y));
    OR4 OR4_291 (.A(OR4_1349_Y), .B(OR4_1014_Y), .C(OR4_1468_Y), .D(
        OR4_1274_Y), .Y(OR4_291_Y));
    OR4 OR4_234 (.A(\R_DATA_TEMPR44[20] ), .B(\R_DATA_TEMPR45[20] ), 
        .C(\R_DATA_TEMPR46[20] ), .D(\R_DATA_TEMPR47[20] ), .Y(
        OR4_234_Y));
    OR4 OR4_1062 (.A(\R_DATA_TEMPR40[13] ), .B(\R_DATA_TEMPR41[13] ), 
        .C(\R_DATA_TEMPR42[13] ), .D(\R_DATA_TEMPR43[13] ), .Y(
        OR4_1062_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%119%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R119C0 (.A_DOUT({
        \R_DATA_TEMPR119[39] , \R_DATA_TEMPR119[38] , 
        \R_DATA_TEMPR119[37] , \R_DATA_TEMPR119[36] , 
        \R_DATA_TEMPR119[35] , \R_DATA_TEMPR119[34] , 
        \R_DATA_TEMPR119[33] , \R_DATA_TEMPR119[32] , 
        \R_DATA_TEMPR119[31] , \R_DATA_TEMPR119[30] , 
        \R_DATA_TEMPR119[29] , \R_DATA_TEMPR119[28] , 
        \R_DATA_TEMPR119[27] , \R_DATA_TEMPR119[26] , 
        \R_DATA_TEMPR119[25] , \R_DATA_TEMPR119[24] , 
        \R_DATA_TEMPR119[23] , \R_DATA_TEMPR119[22] , 
        \R_DATA_TEMPR119[21] , \R_DATA_TEMPR119[20] }), .B_DOUT({
        \R_DATA_TEMPR119[19] , \R_DATA_TEMPR119[18] , 
        \R_DATA_TEMPR119[17] , \R_DATA_TEMPR119[16] , 
        \R_DATA_TEMPR119[15] , \R_DATA_TEMPR119[14] , 
        \R_DATA_TEMPR119[13] , \R_DATA_TEMPR119[12] , 
        \R_DATA_TEMPR119[11] , \R_DATA_TEMPR119[10] , 
        \R_DATA_TEMPR119[9] , \R_DATA_TEMPR119[8] , 
        \R_DATA_TEMPR119[7] , \R_DATA_TEMPR119[6] , 
        \R_DATA_TEMPR119[5] , \R_DATA_TEMPR119[4] , 
        \R_DATA_TEMPR119[3] , \R_DATA_TEMPR119[2] , 
        \R_DATA_TEMPR119[1] , \R_DATA_TEMPR119[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[119][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[29] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[29] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_90 (.A(\R_DATA_TEMPR80[27] ), .B(\R_DATA_TEMPR81[27] ), .C(
        \R_DATA_TEMPR82[27] ), .D(\R_DATA_TEMPR83[27] ), .Y(OR4_90_Y));
    OR4 OR4_1446 (.A(\R_DATA_TEMPR68[7] ), .B(\R_DATA_TEMPR69[7] ), .C(
        \R_DATA_TEMPR70[7] ), .D(\R_DATA_TEMPR71[7] ), .Y(OR4_1446_Y));
    OR4 OR4_1344 (.A(\R_DATA_TEMPR116[10] ), .B(\R_DATA_TEMPR117[10] ), 
        .C(\R_DATA_TEMPR118[10] ), .D(\R_DATA_TEMPR119[10] ), .Y(
        OR4_1344_Y));
    OR4 OR4_46 (.A(\R_DATA_TEMPR112[34] ), .B(\R_DATA_TEMPR113[34] ), 
        .C(\R_DATA_TEMPR114[34] ), .D(\R_DATA_TEMPR115[34] ), .Y(
        OR4_46_Y));
    OR4 OR4_569 (.A(\R_DATA_TEMPR36[4] ), .B(\R_DATA_TEMPR37[4] ), .C(
        \R_DATA_TEMPR38[4] ), .D(\R_DATA_TEMPR39[4] ), .Y(OR4_569_Y));
    OR4 OR4_97 (.A(\R_DATA_TEMPR96[14] ), .B(\R_DATA_TEMPR97[14] ), .C(
        \R_DATA_TEMPR98[14] ), .D(\R_DATA_TEMPR99[14] ), .Y(OR4_97_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%35%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R35C0 (.A_DOUT({
        \R_DATA_TEMPR35[39] , \R_DATA_TEMPR35[38] , 
        \R_DATA_TEMPR35[37] , \R_DATA_TEMPR35[36] , 
        \R_DATA_TEMPR35[35] , \R_DATA_TEMPR35[34] , 
        \R_DATA_TEMPR35[33] , \R_DATA_TEMPR35[32] , 
        \R_DATA_TEMPR35[31] , \R_DATA_TEMPR35[30] , 
        \R_DATA_TEMPR35[29] , \R_DATA_TEMPR35[28] , 
        \R_DATA_TEMPR35[27] , \R_DATA_TEMPR35[26] , 
        \R_DATA_TEMPR35[25] , \R_DATA_TEMPR35[24] , 
        \R_DATA_TEMPR35[23] , \R_DATA_TEMPR35[22] , 
        \R_DATA_TEMPR35[21] , \R_DATA_TEMPR35[20] }), .B_DOUT({
        \R_DATA_TEMPR35[19] , \R_DATA_TEMPR35[18] , 
        \R_DATA_TEMPR35[17] , \R_DATA_TEMPR35[16] , 
        \R_DATA_TEMPR35[15] , \R_DATA_TEMPR35[14] , 
        \R_DATA_TEMPR35[13] , \R_DATA_TEMPR35[12] , 
        \R_DATA_TEMPR35[11] , \R_DATA_TEMPR35[10] , 
        \R_DATA_TEMPR35[9] , \R_DATA_TEMPR35[8] , \R_DATA_TEMPR35[7] , 
        \R_DATA_TEMPR35[6] , \R_DATA_TEMPR35[5] , \R_DATA_TEMPR35[4] , 
        \R_DATA_TEMPR35[3] , \R_DATA_TEMPR35[2] , \R_DATA_TEMPR35[1] , 
        \R_DATA_TEMPR35[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[35][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[8] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[8] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[6]  (.A(OR4_388_Y), .B(OR4_1154_Y), .C(OR4_63_Y), 
        .D(OR4_295_Y), .Y(R_DATA[6]));
    OR4 OR4_592 (.A(\R_DATA_TEMPR12[5] ), .B(\R_DATA_TEMPR13[5] ), .C(
        \R_DATA_TEMPR14[5] ), .D(\R_DATA_TEMPR15[5] ), .Y(OR4_592_Y));
    OR4 OR4_63 (.A(OR4_737_Y), .B(OR4_1036_Y), .C(OR4_502_Y), .D(
        OR4_1357_Y), .Y(OR4_63_Y));
    OR4 OR4_885 (.A(\R_DATA_TEMPR4[7] ), .B(\R_DATA_TEMPR5[7] ), .C(
        \R_DATA_TEMPR6[7] ), .D(\R_DATA_TEMPR7[7] ), .Y(OR4_885_Y));
    OR4 OR4_560 (.A(\R_DATA_TEMPR4[22] ), .B(\R_DATA_TEMPR5[22] ), .C(
        \R_DATA_TEMPR6[22] ), .D(\R_DATA_TEMPR7[22] ), .Y(OR4_560_Y));
    OR4 OR4_217 (.A(\R_DATA_TEMPR8[7] ), .B(\R_DATA_TEMPR9[7] ), .C(
        \R_DATA_TEMPR10[7] ), .D(\R_DATA_TEMPR11[7] ), .Y(OR4_217_Y));
    OR4 OR4_240 (.A(\R_DATA_TEMPR108[10] ), .B(\R_DATA_TEMPR109[10] ), 
        .C(\R_DATA_TEMPR110[10] ), .D(\R_DATA_TEMPR111[10] ), .Y(
        OR4_240_Y));
    OR4 OR4_304 (.A(\R_DATA_TEMPR24[22] ), .B(\R_DATA_TEMPR25[22] ), 
        .C(\R_DATA_TEMPR26[22] ), .D(\R_DATA_TEMPR27[22] ), .Y(
        OR4_304_Y));
    OR4 OR4_117 (.A(OR4_1231_Y), .B(OR4_118_Y), .C(OR4_1257_Y), .D(
        OR4_763_Y), .Y(OR4_117_Y));
    OR4 OR4_1203 (.A(OR4_1241_Y), .B(OR4_747_Y), .C(OR4_728_Y), .D(
        OR4_414_Y), .Y(OR4_1203_Y));
    OR4 OR4_547 (.A(\R_DATA_TEMPR108[11] ), .B(\R_DATA_TEMPR109[11] ), 
        .C(\R_DATA_TEMPR110[11] ), .D(\R_DATA_TEMPR111[11] ), .Y(
        OR4_547_Y));
    OR4 OR4_1413 (.A(\R_DATA_TEMPR48[7] ), .B(\R_DATA_TEMPR49[7] ), .C(
        \R_DATA_TEMPR50[7] ), .D(\R_DATA_TEMPR51[7] ), .Y(OR4_1413_Y));
    OR4 OR4_828 (.A(OR4_57_Y), .B(OR4_548_Y), .C(OR4_520_Y), .D(
        OR4_1300_Y), .Y(OR4_828_Y));
    OR4 OR4_335 (.A(OR4_144_Y), .B(OR4_1528_Y), .C(OR4_1245_Y), .D(
        OR4_51_Y), .Y(OR4_335_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[3]  (.A(CFG3_19_Y), .B(CFG3_2_Y)
        , .Y(\BLKY2[3] ));
    OR4 OR4_1225 (.A(\R_DATA_TEMPR32[24] ), .B(\R_DATA_TEMPR33[24] ), 
        .C(\R_DATA_TEMPR34[24] ), .D(\R_DATA_TEMPR35[24] ), .Y(
        OR4_1225_Y));
    OR4 \OR4_R_DATA[1]  (.A(OR4_1331_Y), .B(OR4_1529_Y), .C(OR4_1077_Y)
        , .D(OR4_866_Y), .Y(R_DATA[1]));
    OR4 OR4_374 (.A(\R_DATA_TEMPR44[37] ), .B(\R_DATA_TEMPR45[37] ), 
        .C(\R_DATA_TEMPR46[37] ), .D(\R_DATA_TEMPR47[37] ), .Y(
        OR4_374_Y));
    OR4 OR4_101 (.A(\R_DATA_TEMPR96[18] ), .B(\R_DATA_TEMPR97[18] ), 
        .C(\R_DATA_TEMPR98[18] ), .D(\R_DATA_TEMPR99[18] ), .Y(
        OR4_101_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[29]  (.A(CFG3_11_Y), .B(
        CFG3_3_Y), .Y(\BLKY2[29] ));
    OR4 OR4_759 (.A(\R_DATA_TEMPR100[29] ), .B(\R_DATA_TEMPR101[29] ), 
        .C(\R_DATA_TEMPR102[29] ), .D(\R_DATA_TEMPR103[29] ), .Y(
        OR4_759_Y));
    OR4 OR4_1521 (.A(\R_DATA_TEMPR8[6] ), .B(\R_DATA_TEMPR9[6] ), .C(
        \R_DATA_TEMPR10[6] ), .D(\R_DATA_TEMPR11[6] ), .Y(OR4_1521_Y));
    OR4 OR4_1636 (.A(\R_DATA_TEMPR56[12] ), .B(\R_DATA_TEMPR57[12] ), 
        .C(\R_DATA_TEMPR58[12] ), .D(\R_DATA_TEMPR59[12] ), .Y(
        OR4_1636_Y));
    OR4 OR4_649 (.A(\R_DATA_TEMPR120[19] ), .B(\R_DATA_TEMPR121[19] ), 
        .C(\R_DATA_TEMPR122[19] ), .D(\R_DATA_TEMPR123[19] ), .Y(
        OR4_649_Y));
    OR4 OR4_594 (.A(\R_DATA_TEMPR8[38] ), .B(\R_DATA_TEMPR9[38] ), .C(
        \R_DATA_TEMPR10[38] ), .D(\R_DATA_TEMPR11[38] ), .Y(OR4_594_Y));
    OR4 OR4_171 (.A(\R_DATA_TEMPR112[11] ), .B(\R_DATA_TEMPR113[11] ), 
        .C(\R_DATA_TEMPR114[11] ), .D(\R_DATA_TEMPR115[11] ), .Y(
        OR4_171_Y));
    OR4 OR4_854 (.A(\R_DATA_TEMPR124[2] ), .B(\R_DATA_TEMPR125[2] ), 
        .C(\R_DATA_TEMPR126[2] ), .D(\R_DATA_TEMPR127[2] ), .Y(
        OR4_854_Y));
    OR4 OR4_1349 (.A(\R_DATA_TEMPR0[33] ), .B(\R_DATA_TEMPR1[33] ), .C(
        \R_DATA_TEMPR2[33] ), .D(\R_DATA_TEMPR3[33] ), .Y(OR4_1349_Y));
    OR4 OR4_713 (.A(OR4_1634_Y), .B(OR2_32_Y), .C(\R_DATA_TEMPR86[34] )
        , .D(\R_DATA_TEMPR87[34] ), .Y(OR4_713_Y));
    OR4 OR4_992 (.A(\R_DATA_TEMPR116[13] ), .B(\R_DATA_TEMPR117[13] ), 
        .C(\R_DATA_TEMPR118[13] ), .D(\R_DATA_TEMPR119[13] ), .Y(
        OR4_992_Y));
    OR4 OR4_553 (.A(OR4_1070_Y), .B(OR4_1396_Y), .C(OR4_830_Y), .D(
        OR4_60_Y), .Y(OR4_553_Y));
    OR4 OR4_1558 (.A(\R_DATA_TEMPR100[2] ), .B(\R_DATA_TEMPR101[2] ), 
        .C(\R_DATA_TEMPR102[2] ), .D(\R_DATA_TEMPR103[2] ), .Y(
        OR4_1558_Y));
    OR4 OR4_1092 (.A(\R_DATA_TEMPR32[9] ), .B(\R_DATA_TEMPR33[9] ), .C(
        \R_DATA_TEMPR34[9] ), .D(\R_DATA_TEMPR35[9] ), .Y(OR4_1092_Y));
    OR4 OR4_1040 (.A(OR4_886_Y), .B(OR4_1183_Y), .C(OR4_637_Y), .D(
        OR4_1500_Y), .Y(OR4_1040_Y));
    OR4 OR4_214 (.A(\R_DATA_TEMPR56[20] ), .B(\R_DATA_TEMPR57[20] ), 
        .C(\R_DATA_TEMPR58[20] ), .D(\R_DATA_TEMPR59[20] ), .Y(
        OR4_214_Y));
    OR4 OR4_246 (.A(\R_DATA_TEMPR92[35] ), .B(\R_DATA_TEMPR93[35] ), 
        .C(\R_DATA_TEMPR94[35] ), .D(\R_DATA_TEMPR95[35] ), .Y(
        OR4_246_Y));
    OR4 OR4_221 (.A(\R_DATA_TEMPR44[13] ), .B(\R_DATA_TEMPR45[13] ), 
        .C(\R_DATA_TEMPR46[13] ), .D(\R_DATA_TEMPR47[13] ), .Y(
        OR4_221_Y));
    OR4 OR4_401 (.A(\R_DATA_TEMPR104[23] ), .B(\R_DATA_TEMPR105[23] ), 
        .C(\R_DATA_TEMPR106[23] ), .D(\R_DATA_TEMPR107[23] ), .Y(
        OR4_401_Y));
    OR4 OR4_1109 (.A(\R_DATA_TEMPR32[14] ), .B(\R_DATA_TEMPR33[14] ), 
        .C(\R_DATA_TEMPR34[14] ), .D(\R_DATA_TEMPR35[14] ), .Y(
        OR4_1109_Y));
    OR4 OR4_74 (.A(\R_DATA_TEMPR72[2] ), .B(\R_DATA_TEMPR73[2] ), .C(
        \R_DATA_TEMPR74[2] ), .D(\R_DATA_TEMPR75[2] ), .Y(OR4_74_Y));
    OR4 OR4_408 (.A(\R_DATA_TEMPR12[29] ), .B(\R_DATA_TEMPR13[29] ), 
        .C(\R_DATA_TEMPR14[29] ), .D(\R_DATA_TEMPR15[29] ), .Y(
        OR4_408_Y));
    OR4 OR4_1283 (.A(\R_DATA_TEMPR40[33] ), .B(\R_DATA_TEMPR41[33] ), 
        .C(\R_DATA_TEMPR42[33] ), .D(\R_DATA_TEMPR43[33] ), .Y(
        OR4_1283_Y));
    OR4 OR4_1259 (.A(OR4_366_Y), .B(OR4_611_Y), .C(OR4_792_Y), .D(
        OR4_564_Y), .Y(OR4_1259_Y));
    OR4 OR4_732 (.A(\R_DATA_TEMPR80[12] ), .B(\R_DATA_TEMPR81[12] ), 
        .C(\R_DATA_TEMPR82[12] ), .D(\R_DATA_TEMPR83[12] ), .Y(
        OR4_732_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%20%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C0 (.A_DOUT({
        \R_DATA_TEMPR20[39] , \R_DATA_TEMPR20[38] , 
        \R_DATA_TEMPR20[37] , \R_DATA_TEMPR20[36] , 
        \R_DATA_TEMPR20[35] , \R_DATA_TEMPR20[34] , 
        \R_DATA_TEMPR20[33] , \R_DATA_TEMPR20[32] , 
        \R_DATA_TEMPR20[31] , \R_DATA_TEMPR20[30] , 
        \R_DATA_TEMPR20[29] , \R_DATA_TEMPR20[28] , 
        \R_DATA_TEMPR20[27] , \R_DATA_TEMPR20[26] , 
        \R_DATA_TEMPR20[25] , \R_DATA_TEMPR20[24] , 
        \R_DATA_TEMPR20[23] , \R_DATA_TEMPR20[22] , 
        \R_DATA_TEMPR20[21] , \R_DATA_TEMPR20[20] }), .B_DOUT({
        \R_DATA_TEMPR20[19] , \R_DATA_TEMPR20[18] , 
        \R_DATA_TEMPR20[17] , \R_DATA_TEMPR20[16] , 
        \R_DATA_TEMPR20[15] , \R_DATA_TEMPR20[14] , 
        \R_DATA_TEMPR20[13] , \R_DATA_TEMPR20[12] , 
        \R_DATA_TEMPR20[11] , \R_DATA_TEMPR20[10] , 
        \R_DATA_TEMPR20[9] , \R_DATA_TEMPR20[8] , \R_DATA_TEMPR20[7] , 
        \R_DATA_TEMPR20[6] , \R_DATA_TEMPR20[5] , \R_DATA_TEMPR20[4] , 
        \R_DATA_TEMPR20[3] , \R_DATA_TEMPR20[2] , \R_DATA_TEMPR20[1] , 
        \R_DATA_TEMPR20[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1563 (.A(OR4_1129_Y), .B(OR4_878_Y), .C(OR4_596_Y), .D(
        OR4_615_Y), .Y(OR4_1563_Y));
    OR4 OR4_471 (.A(\R_DATA_TEMPR60[20] ), .B(\R_DATA_TEMPR61[20] ), 
        .C(\R_DATA_TEMPR62[20] ), .D(\R_DATA_TEMPR63[20] ), .Y(
        OR4_471_Y));
    OR4 OR4_363 (.A(\R_DATA_TEMPR116[17] ), .B(\R_DATA_TEMPR117[17] ), 
        .C(\R_DATA_TEMPR118[17] ), .D(\R_DATA_TEMPR119[17] ), .Y(
        OR4_363_Y));
    OR4 OR4_760 (.A(\R_DATA_TEMPR64[18] ), .B(\R_DATA_TEMPR65[18] ), 
        .C(\R_DATA_TEMPR66[18] ), .D(\R_DATA_TEMPR67[18] ), .Y(
        OR4_760_Y));
    OR4 OR4_391 (.A(\R_DATA_TEMPR8[32] ), .B(\R_DATA_TEMPR9[32] ), .C(
        \R_DATA_TEMPR10[32] ), .D(\R_DATA_TEMPR11[32] ), .Y(OR4_391_Y));
    OR4 OR4_478 (.A(\R_DATA_TEMPR32[1] ), .B(\R_DATA_TEMPR33[1] ), .C(
        \R_DATA_TEMPR34[1] ), .D(\R_DATA_TEMPR35[1] ), .Y(OR4_478_Y));
    OR4 OR4_936 (.A(\R_DATA_TEMPR64[30] ), .B(\R_DATA_TEMPR65[30] ), 
        .C(\R_DATA_TEMPR66[30] ), .D(\R_DATA_TEMPR67[30] ), .Y(
        OR4_936_Y));
    OR4 OR4_644 (.A(\R_DATA_TEMPR8[24] ), .B(\R_DATA_TEMPR9[24] ), .C(
        \R_DATA_TEMPR10[24] ), .D(\R_DATA_TEMPR11[24] ), .Y(OR4_644_Y));
    OR4 OR4_61 (.A(\R_DATA_TEMPR56[31] ), .B(\R_DATA_TEMPR57[31] ), .C(
        \R_DATA_TEMPR58[31] ), .D(\R_DATA_TEMPR59[31] ), .Y(OR4_61_Y));
    OR4 OR4_462 (.A(OR4_1218_Y), .B(OR4_156_Y), .C(OR4_946_Y), .D(
        OR4_1204_Y), .Y(OR4_462_Y));
    OR4 OR4_1034 (.A(\R_DATA_TEMPR8[39] ), .B(\R_DATA_TEMPR9[39] ), .C(
        \R_DATA_TEMPR10[39] ), .D(\R_DATA_TEMPR11[39] ), .Y(OR4_1034_Y)
        );
    OR4 OR4_1449 (.A(\R_DATA_TEMPR48[1] ), .B(\R_DATA_TEMPR49[1] ), .C(
        \R_DATA_TEMPR50[1] ), .D(\R_DATA_TEMPR51[1] ), .Y(OR4_1449_Y));
    OR4 OR4_635 (.A(\R_DATA_TEMPR72[6] ), .B(\R_DATA_TEMPR73[6] ), .C(
        \R_DATA_TEMPR74[6] ), .D(\R_DATA_TEMPR75[6] ), .Y(OR4_635_Y));
    OR4 OR4_522 (.A(\R_DATA_TEMPR112[17] ), .B(\R_DATA_TEMPR113[17] ), 
        .C(\R_DATA_TEMPR114[17] ), .D(\R_DATA_TEMPR115[17] ), .Y(
        OR4_522_Y));
    OR4 OR4_686 (.A(\R_DATA_TEMPR4[14] ), .B(\R_DATA_TEMPR5[14] ), .C(
        \R_DATA_TEMPR6[14] ), .D(\R_DATA_TEMPR7[14] ), .Y(OR4_686_Y));
    OR2 OR2_5 (.A(\R_DATA_TEMPR84[39] ), .B(\R_DATA_TEMPR85[39] ), .Y(
        OR2_5_Y));
    OR4 OR4_315 (.A(\R_DATA_TEMPR124[32] ), .B(\R_DATA_TEMPR125[32] ), 
        .C(\R_DATA_TEMPR126[32] ), .D(\R_DATA_TEMPR127[32] ), .Y(
        OR4_315_Y));
    OR4 OR4_469 (.A(\R_DATA_TEMPR60[2] ), .B(\R_DATA_TEMPR61[2] ), .C(
        \R_DATA_TEMPR62[2] ), .D(\R_DATA_TEMPR63[2] ), .Y(OR4_469_Y));
    OR4 OR4_1333 (.A(\R_DATA_TEMPR32[36] ), .B(\R_DATA_TEMPR33[36] ), 
        .C(\R_DATA_TEMPR34[36] ), .D(\R_DATA_TEMPR35[36] ), .Y(
        OR4_1333_Y));
    OR4 OR4_490 (.A(\R_DATA_TEMPR88[14] ), .B(\R_DATA_TEMPR89[14] ), 
        .C(\R_DATA_TEMPR90[14] ), .D(\R_DATA_TEMPR91[14] ), .Y(
        OR4_490_Y));
    OR4 OR4_40 (.A(\R_DATA_TEMPR12[8] ), .B(\R_DATA_TEMPR13[8] ), .C(
        \R_DATA_TEMPR14[8] ), .D(\R_DATA_TEMPR15[8] ), .Y(OR4_40_Y));
    OR4 OR4_509 (.A(\R_DATA_TEMPR20[6] ), .B(\R_DATA_TEMPR21[6] ), .C(
        \R_DATA_TEMPR22[6] ), .D(\R_DATA_TEMPR23[6] ), .Y(OR4_509_Y));
    OR4 OR4_166 (.A(\R_DATA_TEMPR108[29] ), .B(\R_DATA_TEMPR109[29] ), 
        .C(\R_DATA_TEMPR110[29] ), .D(\R_DATA_TEMPR111[29] ), .Y(
        OR4_166_Y));
    OR4 OR4_1189 (.A(\R_DATA_TEMPR20[35] ), .B(\R_DATA_TEMPR21[35] ), 
        .C(\R_DATA_TEMPR22[35] ), .D(\R_DATA_TEMPR23[35] ), .Y(
        OR4_1189_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[26]  (.A(CFG3_0_Y), .B(CFG3_3_Y)
        , .Y(\BLKY2[26] ));
    OR4 OR4_500 (.A(\R_DATA_TEMPR0[5] ), .B(\R_DATA_TEMPR1[5] ), .C(
        \R_DATA_TEMPR2[5] ), .D(\R_DATA_TEMPR3[5] ), .Y(OR4_500_Y));
    OR4 OR4_1574 (.A(OR4_182_Y), .B(OR4_820_Y), .C(OR4_1366_Y), .D(
        OR4_753_Y), .Y(OR4_1574_Y));
    OR4 OR4_47 (.A(OR4_685_Y), .B(OR4_997_Y), .C(OR4_1247_Y), .D(
        OR4_1046_Y), .Y(OR4_47_Y));
    OR4 OR4_1626 (.A(\R_DATA_TEMPR12[12] ), .B(\R_DATA_TEMPR13[12] ), 
        .C(\R_DATA_TEMPR14[12] ), .D(\R_DATA_TEMPR15[12] ), .Y(
        OR4_1626_Y));
    OR4 OR4_1106 (.A(OR4_347_Y), .B(OR2_27_Y), .C(\R_DATA_TEMPR86[19] )
        , .D(\R_DATA_TEMPR87[19] ), .Y(OR4_1106_Y));
    OR4 OR4_579 (.A(\R_DATA_TEMPR28[13] ), .B(\R_DATA_TEMPR29[13] ), 
        .C(\R_DATA_TEMPR30[13] ), .D(\R_DATA_TEMPR31[13] ), .Y(
        OR4_579_Y));
    OR4 OR4_1113 (.A(\R_DATA_TEMPR68[28] ), .B(\R_DATA_TEMPR69[28] ), 
        .C(\R_DATA_TEMPR70[28] ), .D(\R_DATA_TEMPR71[28] ), .Y(
        OR4_1113_Y));
    OR4 OR4_1401 (.A(\R_DATA_TEMPR76[5] ), .B(\R_DATA_TEMPR77[5] ), .C(
        \R_DATA_TEMPR78[5] ), .D(\R_DATA_TEMPR79[5] ), .Y(OR4_1401_Y));
    OR4 OR4_570 (.A(\R_DATA_TEMPR76[21] ), .B(\R_DATA_TEMPR77[21] ), 
        .C(\R_DATA_TEMPR78[21] ), .D(\R_DATA_TEMPR79[21] ), .Y(
        OR4_570_Y));
    OR4 OR4_1375 (.A(\R_DATA_TEMPR124[35] ), .B(\R_DATA_TEMPR125[35] ), 
        .C(\R_DATA_TEMPR126[35] ), .D(\R_DATA_TEMPR127[35] ), .Y(
        OR4_1375_Y));
    OR4 OR4_524 (.A(\R_DATA_TEMPR104[15] ), .B(\R_DATA_TEMPR105[15] ), 
        .C(\R_DATA_TEMPR106[15] ), .D(\R_DATA_TEMPR107[15] ), .Y(
        OR4_524_Y));
    OR4 OR4_1201 (.A(\R_DATA_TEMPR68[15] ), .B(\R_DATA_TEMPR69[15] ), 
        .C(\R_DATA_TEMPR70[15] ), .D(\R_DATA_TEMPR71[15] ), .Y(
        OR4_1201_Y));
    OR4 OR4_1108 (.A(\R_DATA_TEMPR68[3] ), .B(\R_DATA_TEMPR69[3] ), .C(
        \R_DATA_TEMPR70[3] ), .D(\R_DATA_TEMPR71[3] ), .Y(OR4_1108_Y));
    OR4 \OR4_R_DATA[28]  (.A(OR4_1431_Y), .B(OR4_1198_Y), .C(OR4_462_Y)
        , .D(OR4_679_Y), .Y(R_DATA[28]));
    RAM1K20 #( .RAMINDEX("PF_SRAM%65536-65536%40-40%POWER%11%0%TWO-PORT%ECC_EN-0")
         )  PF_SRAM_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C0 (.A_DOUT({
        \R_DATA_TEMPR11[39] , \R_DATA_TEMPR11[38] , 
        \R_DATA_TEMPR11[37] , \R_DATA_TEMPR11[36] , 
        \R_DATA_TEMPR11[35] , \R_DATA_TEMPR11[34] , 
        \R_DATA_TEMPR11[33] , \R_DATA_TEMPR11[32] , 
        \R_DATA_TEMPR11[31] , \R_DATA_TEMPR11[30] , 
        \R_DATA_TEMPR11[29] , \R_DATA_TEMPR11[28] , 
        \R_DATA_TEMPR11[27] , \R_DATA_TEMPR11[26] , 
        \R_DATA_TEMPR11[25] , \R_DATA_TEMPR11[24] , 
        \R_DATA_TEMPR11[23] , \R_DATA_TEMPR11[22] , 
        \R_DATA_TEMPR11[21] , \R_DATA_TEMPR11[20] }), .B_DOUT({
        \R_DATA_TEMPR11[19] , \R_DATA_TEMPR11[18] , 
        \R_DATA_TEMPR11[17] , \R_DATA_TEMPR11[16] , 
        \R_DATA_TEMPR11[15] , \R_DATA_TEMPR11[14] , 
        \R_DATA_TEMPR11[13] , \R_DATA_TEMPR11[12] , 
        \R_DATA_TEMPR11[11] , \R_DATA_TEMPR11[10] , 
        \R_DATA_TEMPR11[9] , \R_DATA_TEMPR11[8] , \R_DATA_TEMPR11[7] , 
        \R_DATA_TEMPR11[6] , \R_DATA_TEMPR11[5] , \R_DATA_TEMPR11[4] , 
        \R_DATA_TEMPR11[3] , \R_DATA_TEMPR11[2] , \R_DATA_TEMPR11[1] , 
        \R_DATA_TEMPR11[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[2] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_922 (.A(OR4_1031_Y), .B(OR4_1306_Y), .C(OR4_802_Y), .D(
        OR4_552_Y), .Y(OR4_922_Y));
    OR4 OR4_368 (.A(\R_DATA_TEMPR100[1] ), .B(\R_DATA_TEMPR101[1] ), 
        .C(\R_DATA_TEMPR102[1] ), .D(\R_DATA_TEMPR103[1] ), .Y(
        OR4_368_Y));
    OR4 OR4_1593 (.A(\R_DATA_TEMPR4[37] ), .B(\R_DATA_TEMPR5[37] ), .C(
        \R_DATA_TEMPR6[37] ), .D(\R_DATA_TEMPR7[37] ), .Y(OR4_1593_Y));
    OR4 OR4_1519 (.A(\R_DATA_TEMPR68[2] ), .B(\R_DATA_TEMPR69[2] ), .C(
        \R_DATA_TEMPR70[2] ), .D(\R_DATA_TEMPR71[2] ), .Y(OR4_1519_Y));
    OR4 OR4_712 (.A(\R_DATA_TEMPR112[28] ), .B(\R_DATA_TEMPR113[28] ), 
        .C(\R_DATA_TEMPR114[28] ), .D(\R_DATA_TEMPR115[28] ), .Y(
        OR4_712_Y));
    OR4 OR4_630 (.A(\R_DATA_TEMPR108[31] ), .B(\R_DATA_TEMPR109[31] ), 
        .C(\R_DATA_TEMPR110[31] ), .D(\R_DATA_TEMPR111[31] ), .Y(
        OR4_630_Y));
    OR4 OR4_916 (.A(\R_DATA_TEMPR40[34] ), .B(\R_DATA_TEMPR41[34] ), 
        .C(\R_DATA_TEMPR42[34] ), .D(\R_DATA_TEMPR43[34] ), .Y(
        OR4_916_Y));
    OR4 OR4_98 (.A(\R_DATA_TEMPR124[12] ), .B(\R_DATA_TEMPR125[12] ), 
        .C(\R_DATA_TEMPR126[12] ), .D(\R_DATA_TEMPR127[12] ), .Y(
        OR4_98_Y));
    OR4 OR4_1024 (.A(\R_DATA_TEMPR104[21] ), .B(\R_DATA_TEMPR105[21] ), 
        .C(\R_DATA_TEMPR106[21] ), .D(\R_DATA_TEMPR107[21] ), .Y(
        OR4_1024_Y));
    OR4 OR4_321 (.A(OR4_296_Y), .B(OR2_21_Y), .C(\R_DATA_TEMPR86[5] ), 
        .D(\R_DATA_TEMPR87[5] ), .Y(OR4_321_Y));
    OR4 OR4_1186 (.A(\R_DATA_TEMPR16[29] ), .B(\R_DATA_TEMPR17[29] ), 
        .C(\R_DATA_TEMPR18[29] ), .D(\R_DATA_TEMPR19[29] ), .Y(
        OR4_1186_Y));
    OR4 OR4_615 (.A(\R_DATA_TEMPR124[27] ), .B(\R_DATA_TEMPR125[27] ), 
        .C(\R_DATA_TEMPR126[27] ), .D(\R_DATA_TEMPR127[27] ), .Y(
        OR4_615_Y));
    OR4 OR4_1481 (.A(\R_DATA_TEMPR12[14] ), .B(\R_DATA_TEMPR13[14] ), 
        .C(\R_DATA_TEMPR14[14] ), .D(\R_DATA_TEMPR15[14] ), .Y(
        OR4_1481_Y));
    OR4 OR4_1440 (.A(\R_DATA_TEMPR120[22] ), .B(\R_DATA_TEMPR121[22] ), 
        .C(\R_DATA_TEMPR122[22] ), .D(\R_DATA_TEMPR123[22] ), .Y(
        OR4_1440_Y));
    OR4 OR4_337 (.A(\R_DATA_TEMPR108[15] ), .B(\R_DATA_TEMPR109[15] ), 
        .C(\R_DATA_TEMPR110[15] ), .D(\R_DATA_TEMPR111[15] ), .Y(
        OR4_337_Y));
    OR4 OR4_130 (.A(OR4_1310_Y), .B(OR4_1027_Y), .C(OR4_752_Y), .D(
        OR4_1573_Y), .Y(OR4_130_Y));
    OR2 OR2_25 (.A(\R_DATA_TEMPR84[33] ), .B(\R_DATA_TEMPR85[33] ), .Y(
        OR2_25_Y));
    OR4 OR4_1323 (.A(OR4_810_Y), .B(OR4_681_Y), .C(OR4_1224_Y), .D(
        OR4_619_Y), .Y(OR4_1323_Y));
    OR4 OR4_1036 (.A(\R_DATA_TEMPR100[6] ), .B(\R_DATA_TEMPR101[6] ), 
        .C(\R_DATA_TEMPR102[6] ), .D(\R_DATA_TEMPR103[6] ), .Y(
        OR4_1036_Y));
    OR4 OR4_1281 (.A(\R_DATA_TEMPR80[4] ), .B(\R_DATA_TEMPR81[4] ), .C(
        \R_DATA_TEMPR82[4] ), .D(\R_DATA_TEMPR83[4] ), .Y(OR4_1281_Y));
    OR4 OR4_169 (.A(\R_DATA_TEMPR48[23] ), .B(\R_DATA_TEMPR49[23] ), 
        .C(\R_DATA_TEMPR50[23] ), .D(\R_DATA_TEMPR51[23] ), .Y(
        OR4_169_Y));
    OR4 OR4_303 (.A(\R_DATA_TEMPR72[29] ), .B(\R_DATA_TEMPR73[29] ), 
        .C(\R_DATA_TEMPR74[29] ), .D(\R_DATA_TEMPR75[29] ), .Y(
        OR4_303_Y));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
