///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: MUX_DDR_simulator.v
// File history:
//      <v1.0: <04/2021>: First version
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// MUX DTC Data Request signals from Top_Serde to use DDR simulator pattern.
// N.B.: Only pattern = 0 (increasing counter) is generated by DDR simulator.
//
// Targeted device: <Family::PolarFire> <Die::MPF300TS> <Package::FCG1152>
// Author: Monica Tecchio
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

//`timescale <time_units> / <precision>

module MUX_DDR_simulator( 
	input					RDOUT_CLK,
   input					DDRSIM_EN,  // if 0, DDR packets to Top_Serdes;  if 1, DDR_Simulator packets to Top_Serdes
   input					DDR_DDR3_FULL,
   input					DDR_DATA_READY,
   input					DDR_LAST_WORD,
   input    [31:0]	DDR_WR_CNT,
   input    [31:0]	DDR_RD_CNT,
   input    [31:0]	DDR_FIFO_RD_CNT,
   input    [15:0]	DDR_DATA_PCKTS,
   input    [63:0]   DDR_DATA,
   input					DDRSIM_DDR3_FULL,
   input					DDRSIM_DATA_READY,
   input					DDRSIM_LAST_WORD,
   input    [31:0]	DDRSIM_WR_CNT,
   input    [31:0]	DDRSIM_RD_CNT,
   input    [31:0]	DDRSIM_FIFO_RD_CNT,
   input    [15:0]	DDRSIM_DATA_PCKTS,
   input    [63:0]   DDRSIM_DATA,
	output reg			DDR3_FULL,
	output reg			MEMFIFO_DATA_READY,
	output reg			MEMFIFO_LAST_WORD,
   output reg [31:0]	MEM_WR_CNT,
   output reg [31:0]	MEM_RD_CNT,
   output reg [31:0]	MEMFIFO_RD_CNT,
   output reg [15:0]	MEMFIFO_DATA_PCKTS,
   output reg [63:0]	MEMFIFO_DATA
  );

   always @ (*)
   begin
		DDR3_FULL 	   	= (DDRSIM_EN==1'b1) ? DDRSIM_DDR3_FULL  	: DDR_DDR3_FULL;
		MEMFIFO_DATA_READY= (DDRSIM_EN==1'b1) ? DDRSIM_DATA_READY 	: DDR_DATA_READY;
		MEMFIFO_LAST_WORD	= (DDRSIM_EN==1'b1) ? DDRSIM_LAST_WORD  	: DDR_LAST_WORD;
		MEM_WR_CNT			= (DDRSIM_EN==1'b1) ? DDRSIM_WR_CNT			: DDR_WR_CNT;
		MEM_RD_CNT			= (DDRSIM_EN==1'b1) ? DDRSIM_RD_CNT			: DDR_RD_CNT;
		MEMFIFO_RD_CNT		= (DDRSIM_EN==1'b1) ? DDRSIM_FIFO_RD_CNT	: DDR_FIFO_RD_CNT;
		MEMFIFO_DATA_PCKTS= (DDRSIM_EN==1'b1) ? DDRSIM_DATA_PCKTS	: DDR_DATA_PCKTS;
		MEMFIFO_DATA		= (DDRSIM_EN==1'b1) ? DDRSIM_DATA			: DDR_DATA;
  end

  
endmodule

